module FFT1024_LUT(n, twiddle);
	input [9:0] n;
		
	output reg [31:0] twiddle;
	
	always @ (n)
	begin
		//$display("LUT address=%d", n);
		case(n)
		10'd0  : twiddle = { 16'd32767   ,  16'd0       }; //i=0  n=1024 twiddle= 1               + i 0
		10'd1  : twiddle = { 16'd32766   , -16'd201     }; //i=1  n=1024 twiddle= 9.999812e-01    + i -6.135885e-03
		10'd2  : twiddle = { 16'd32765   , -16'd402     }; //i=2  n=1024 twiddle= 9.999247e-01    + i -1.227154e-02
		10'd3  : twiddle = { 16'd32761   , -16'd603     }; //i=3  n=1024 twiddle= 9.998306e-01    + i -1.840673e-02
		10'd4  : twiddle = { 16'd32757   , -16'd804     }; //i=4  n=1024 twiddle= 9.996988e-01    + i -2.454123e-02
		10'd5  : twiddle = { 16'd32752   , -16'd1005    }; //i=5  n=1024 twiddle= 9.995294e-01    + i -3.067480e-02
		10'd6  : twiddle = { 16'd32745   , -16'd1206    }; //i=6  n=1024 twiddle= 9.993224e-01    + i -3.680722e-02
		10'd7  : twiddle = { 16'd32737   , -16'd1407    }; //i=7  n=1024 twiddle= 9.990777e-01    + i -4.293826e-02
		10'd8  : twiddle = { 16'd32728   , -16'd1608    }; //i=8  n=1024 twiddle= 9.987955e-01    + i -4.906767e-02
		10'd9  : twiddle = { 16'd32717   , -16'd1809    }; //i=9  n=1024 twiddle= 9.984756e-01    + i -5.519524e-02
		10'd10 : twiddle = { 16'd32705   , -16'd2009    }; //i=10 n=1024 twiddle= 9.981181e-01    + i -6.132074e-02
		10'd11 : twiddle = { 16'd32692   , -16'd2210    }; //i=11 n=1024 twiddle= 9.977231e-01    + i -6.744392e-02
		10'd12 : twiddle = { 16'd32678   , -16'd2410    }; //i=12 n=1024 twiddle= 9.972905e-01    + i -7.356456e-02
		10'd13 : twiddle = { 16'd32663   , -16'd2611    }; //i=13 n=1024 twiddle= 9.968203e-01    + i -7.968244e-02
		10'd14 : twiddle = { 16'd32646   , -16'd2811    }; //i=14 n=1024 twiddle= 9.963126e-01    + i -8.579731e-02
		10'd15 : twiddle = { 16'd32628   , -16'd3012    }; //i=15 n=1024 twiddle= 9.957674e-01    + i -9.190896e-02
		10'd16 : twiddle = { 16'd32609   , -16'd3212    }; //i=16 n=1024 twiddle= 9.951847e-01    + i -9.801714e-02
		10'd17 : twiddle = { 16'd32589   , -16'd3412    }; //i=17 n=1024 twiddle= 9.945646e-01    + i -1.041216e-01
		10'd18 : twiddle = { 16'd32567   , -16'd3612    }; //i=18 n=1024 twiddle= 9.939070e-01    + i -1.102222e-01
		10'd19 : twiddle = { 16'd32545   , -16'd3811    }; //i=19 n=1024 twiddle= 9.932119e-01    + i -1.163186e-01
		10'd20 : twiddle = { 16'd32521   , -16'd4011    }; //i=20 n=1024 twiddle= 9.924795e-01    + i -1.224107e-01
		10'd21 : twiddle = { 16'd32495   , -16'd4210    }; //i=21 n=1024 twiddle= 9.917098e-01    + i -1.284981e-01
		10'd22 : twiddle = { 16'd32469   , -16'd4410    }; //i=22 n=1024 twiddle= 9.909026e-01    + i -1.345807e-01
		10'd23 : twiddle = { 16'd32441   , -16'd4609    }; //i=23 n=1024 twiddle= 9.900582e-01    + i -1.406582e-01
		10'd24 : twiddle = { 16'd32412   , -16'd4808    }; //i=24 n=1024 twiddle= 9.891765e-01    + i -1.467305e-01
		10'd25 : twiddle = { 16'd32382   , -16'd5007    }; //i=25 n=1024 twiddle= 9.882576e-01    + i -1.527972e-01
		10'd26 : twiddle = { 16'd32351   , -16'd5205    }; //i=26 n=1024 twiddle= 9.873014e-01    + i -1.588581e-01
		10'd27 : twiddle = { 16'd32318   , -16'd5404    }; //i=27 n=1024 twiddle= 9.863081e-01    + i -1.649131e-01
		10'd28 : twiddle = { 16'd32285   , -16'd5602    }; //i=28 n=1024 twiddle= 9.852776e-01    + i -1.709619e-01
		10'd29 : twiddle = { 16'd32250   , -16'd5800    }; //i=29 n=1024 twiddle= 9.842101e-01    + i -1.770042e-01
		10'd30 : twiddle = { 16'd32213   , -16'd5998    }; //i=30 n=1024 twiddle= 9.831055e-01    + i -1.830399e-01
		10'd31 : twiddle = { 16'd32176   , -16'd6195    }; //i=31 n=1024 twiddle= 9.819639e-01    + i -1.890687e-01
		10'd32 : twiddle = { 16'd32137   , -16'd6393    }; //i=32 n=1024 twiddle= 9.807853e-01    + i -1.950903e-01
		10'd33 : twiddle = { 16'd32098   , -16'd6590    }; //i=33 n=1024 twiddle= 9.795698e-01    + i -2.011046e-01
		10'd34 : twiddle = { 16'd32057   , -16'd6786    }; //i=34 n=1024 twiddle= 9.783174e-01    + i -2.071114e-01
		10'd35 : twiddle = { 16'd32014   , -16'd6983    }; //i=35 n=1024 twiddle= 9.770281e-01    + i -2.131103e-01
		10'd36 : twiddle = { 16'd31971   , -16'd7179    }; //i=36 n=1024 twiddle= 9.757021e-01    + i -2.191012e-01
		10'd37 : twiddle = { 16'd31926   , -16'd7375    }; //i=37 n=1024 twiddle= 9.743394e-01    + i -2.250839e-01
		10'd38 : twiddle = { 16'd31880   , -16'd7571    }; //i=38 n=1024 twiddle= 9.729400e-01    + i -2.310581e-01
		10'd39 : twiddle = { 16'd31833   , -16'd7767    }; //i=39 n=1024 twiddle= 9.715039e-01    + i -2.370236e-01
		10'd40 : twiddle = { 16'd31785   , -16'd7962    }; //i=40 n=1024 twiddle= 9.700313e-01    + i -2.429802e-01
		10'd41 : twiddle = { 16'd31736   , -16'd8157    }; //i=41 n=1024 twiddle= 9.685221e-01    + i -2.489276e-01
		10'd42 : twiddle = { 16'd31685   , -16'd8351    }; //i=42 n=1024 twiddle= 9.669765e-01    + i -2.548657e-01
		10'd43 : twiddle = { 16'd31633   , -16'd8545    }; //i=43 n=1024 twiddle= 9.653944e-01    + i -2.607941e-01
		10'd44 : twiddle = { 16'd31580   , -16'd8739    }; //i=44 n=1024 twiddle= 9.637761e-01    + i -2.667128e-01
		10'd45 : twiddle = { 16'd31526   , -16'd8933    }; //i=45 n=1024 twiddle= 9.621214e-01    + i -2.726214e-01
		10'd46 : twiddle = { 16'd31470   , -16'd9126    }; //i=46 n=1024 twiddle= 9.604305e-01    + i -2.785197e-01
		10'd47 : twiddle = { 16'd31414   , -16'd9319    }; //i=47 n=1024 twiddle= 9.587035e-01    + i -2.844075e-01
		10'd48 : twiddle = { 16'd31356   , -16'd9512    }; //i=48 n=1024 twiddle= 9.569403e-01    + i -2.902847e-01
		10'd49 : twiddle = { 16'd31297   , -16'd9704    }; //i=49 n=1024 twiddle= 9.551412e-01    + i -2.961509e-01
		10'd50 : twiddle = { 16'd31237   , -16'd9896    }; //i=50 n=1024 twiddle= 9.533060e-01    + i -3.020059e-01
		10'd51 : twiddle = { 16'd31176   , -16'd10087   }; //i=51 n=1024 twiddle= 9.514350e-01    + i -3.078496e-01
		10'd52 : twiddle = { 16'd31113   , -16'd10278   }; //i=52 n=1024 twiddle= 9.495282e-01    + i -3.136817e-01
		10'd53 : twiddle = { 16'd31050   , -16'd10469   }; //i=53 n=1024 twiddle= 9.475856e-01    + i -3.195020e-01
		10'd54 : twiddle = { 16'd30985   , -16'd10659   }; //i=54 n=1024 twiddle= 9.456073e-01    + i -3.253103e-01
		10'd55 : twiddle = { 16'd30919   , -16'd10849   }; //i=55 n=1024 twiddle= 9.435935e-01    + i -3.311063e-01
		10'd56 : twiddle = { 16'd30852   , -16'd11039   }; //i=56 n=1024 twiddle= 9.415441e-01    + i -3.368899e-01
		10'd57 : twiddle = { 16'd30783   , -16'd11228   }; //i=57 n=1024 twiddle= 9.394592e-01    + i -3.426607e-01
		10'd58 : twiddle = { 16'd30714   , -16'd11417   }; //i=58 n=1024 twiddle= 9.373390e-01    + i -3.484187e-01
		10'd59 : twiddle = { 16'd30643   , -16'd11605   }; //i=59 n=1024 twiddle= 9.351835e-01    + i -3.541635e-01
		10'd60 : twiddle = { 16'd30571   , -16'd11793   }; //i=60 n=1024 twiddle= 9.329928e-01    + i -3.598950e-01
		10'd61 : twiddle = { 16'd30498   , -16'd11980   }; //i=61 n=1024 twiddle= 9.307670e-01    + i -3.656130e-01
		10'd62 : twiddle = { 16'd30424   , -16'd12167   }; //i=62 n=1024 twiddle= 9.285061e-01    + i -3.713172e-01
		10'd63 : twiddle = { 16'd30349   , -16'd12353   }; //i=63 n=1024 twiddle= 9.262102e-01    + i -3.770074e-01
		10'd64 : twiddle = { 16'd30273   , -16'd12539   }; //i=64 n=1024 twiddle= 9.238795e-01    + i -3.826834e-01
		10'd65 : twiddle = { 16'd30195   , -16'd12725   }; //i=65 n=1024 twiddle= 9.215140e-01    + i -3.883450e-01
		10'd66 : twiddle = { 16'd30117   , -16'd12910   }; //i=66 n=1024 twiddle= 9.191139e-01    + i -3.939920e-01
		10'd67 : twiddle = { 16'd30037   , -16'd13094   }; //i=67 n=1024 twiddle= 9.166791e-01    + i -3.996242e-01
		10'd68 : twiddle = { 16'd29956   , -16'd13279   }; //i=68 n=1024 twiddle= 9.142098e-01    + i -4.052413e-01
		10'd69 : twiddle = { 16'd29874   , -16'd13462   }; //i=69 n=1024 twiddle= 9.117060e-01    + i -4.108432e-01
		10'd70 : twiddle = { 16'd29791   , -16'd13645   }; //i=70 n=1024 twiddle= 9.091680e-01    + i -4.164296e-01
		10'd71 : twiddle = { 16'd29706   , -16'd13828   }; //i=71 n=1024 twiddle= 9.065957e-01    + i -4.220003e-01
		10'd72 : twiddle = { 16'd29621   , -16'd14010   }; //i=72 n=1024 twiddle= 9.039893e-01    + i -4.275551e-01
		10'd73 : twiddle = { 16'd29534   , -16'd14191   }; //i=73 n=1024 twiddle= 9.013488e-01    + i -4.330938e-01
		10'd74 : twiddle = { 16'd29447   , -16'd14372   }; //i=74 n=1024 twiddle= 8.986745e-01    + i -4.386162e-01
		10'd75 : twiddle = { 16'd29358   , -16'd14553   }; //i=75 n=1024 twiddle= 8.959662e-01    + i -4.441221e-01
		10'd76 : twiddle = { 16'd29268   , -16'd14732   }; //i=76 n=1024 twiddle= 8.932243e-01    + i -4.496113e-01
		10'd77 : twiddle = { 16'd29177   , -16'd14912   }; //i=77 n=1024 twiddle= 8.904487e-01    + i -4.550836e-01
		10'd78 : twiddle = { 16'd29085   , -16'd15090   }; //i=78 n=1024 twiddle= 8.876396e-01    + i -4.605387e-01
		10'd79 : twiddle = { 16'd28992   , -16'd15269   }; //i=79 n=1024 twiddle= 8.847971e-01    + i -4.659765e-01
		10'd80 : twiddle = { 16'd28898   , -16'd15446   }; //i=80 n=1024 twiddle= 8.819213e-01    + i -4.713967e-01
		10'd81 : twiddle = { 16'd28803   , -16'd15623   }; //i=81 n=1024 twiddle= 8.790122e-01    + i -4.767992e-01
		10'd82 : twiddle = { 16'd28706   , -16'd15800   }; //i=82 n=1024 twiddle= 8.760701e-01    + i -4.821838e-01
		10'd83 : twiddle = { 16'd28609   , -16'd15976   }; //i=83 n=1024 twiddle= 8.730950e-01    + i -4.875502e-01
		10'd84 : twiddle = { 16'd28510   , -16'd16151   }; //i=84 n=1024 twiddle= 8.700870e-01    + i -4.928982e-01
		10'd85 : twiddle = { 16'd28411   , -16'd16325   }; //i=85 n=1024 twiddle= 8.670462e-01    + i -4.982277e-01
		10'd86 : twiddle = { 16'd28310   , -16'd16499   }; //i=86 n=1024 twiddle= 8.639729e-01    + i -5.035384e-01
		10'd87 : twiddle = { 16'd28208   , -16'd16673   }; //i=87 n=1024 twiddle= 8.608669e-01    + i -5.088301e-01
		10'd88 : twiddle = { 16'd28105   , -16'd16846   }; //i=88 n=1024 twiddle= 8.577286e-01    + i -5.141027e-01
		10'd89 : twiddle = { 16'd28001   , -16'd17018   }; //i=89 n=1024 twiddle= 8.545580e-01    + i -5.193560e-01
		10'd90 : twiddle = { 16'd27896   , -16'd17189   }; //i=90 n=1024 twiddle= 8.513552e-01    + i -5.245897e-01
		10'd91 : twiddle = { 16'd27790   , -16'd17360   }; //i=91 n=1024 twiddle= 8.481203e-01    + i -5.298036e-01
		10'd92 : twiddle = { 16'd27683   , -16'd17530   }; //i=92 n=1024 twiddle= 8.448536e-01    + i -5.349976e-01
		10'd93 : twiddle = { 16'd27575   , -16'd17700   }; //i=93 n=1024 twiddle= 8.415550e-01    + i -5.401715e-01
		10'd94 : twiddle = { 16'd27466   , -16'd17869   }; //i=94 n=1024 twiddle= 8.382247e-01    + i -5.453250e-01
		10'd95 : twiddle = { 16'd27356   , -16'd18037   }; //i=95 n=1024 twiddle= 8.348629e-01    + i -5.504580e-01
		10'd96 : twiddle = { 16'd27245   , -16'd18204   }; //i=96 n=1024 twiddle= 8.314696e-01    + i -5.555702e-01
		10'd97 : twiddle = { 16'd27133   , -16'd18371   }; //i=97 n=1024 twiddle= 8.280450e-01    + i -5.606616e-01
		10'd98 : twiddle = { 16'd27019   , -16'd18537   }; //i=98 n=1024 twiddle= 8.245893e-01    + i -5.657318e-01
		10'd99 : twiddle = { 16'd26905   , -16'd18703   }; //i=99 n=1024 twiddle= 8.211025e-01    + i -5.707807e-01
		10'd100: twiddle = { 16'd26790   , -16'd18868   }; //i=100 n=1024 twiddle= 8.175848e-01    + i -5.758082e-01
		10'd101: twiddle = { 16'd26674   , -16'd19032   }; //i=101 n=1024 twiddle= 8.140363e-01    + i -5.808140e-01
		10'd102: twiddle = { 16'd26556   , -16'd19195   }; //i=102 n=1024 twiddle= 8.104572e-01    + i -5.857979e-01
		10'd103: twiddle = { 16'd26438   , -16'd19357   }; //i=103 n=1024 twiddle= 8.068476e-01    + i -5.907597e-01
		10'd104: twiddle = { 16'd26319   , -16'd19519   }; //i=104 n=1024 twiddle= 8.032075e-01    + i -5.956993e-01
		10'd105: twiddle = { 16'd26198   , -16'd19680   }; //i=105 n=1024 twiddle= 7.995373e-01    + i -6.006165e-01
		10'd106: twiddle = { 16'd26077   , -16'd19841   }; //i=106 n=1024 twiddle= 7.958369e-01    + i -6.055110e-01
		10'd107: twiddle = { 16'd25955   , -16'd20000   }; //i=107 n=1024 twiddle= 7.921066e-01    + i -6.103828e-01
		10'd108: twiddle = { 16'd25832   , -16'd20159   }; //i=108 n=1024 twiddle= 7.883464e-01    + i -6.152316e-01
		10'd109: twiddle = { 16'd25708   , -16'd20317   }; //i=109 n=1024 twiddle= 7.845566e-01    + i -6.200572e-01
		10'd110: twiddle = { 16'd25582   , -16'd20475   }; //i=110 n=1024 twiddle= 7.807372e-01    + i -6.248595e-01
		10'd111: twiddle = { 16'd25456   , -16'd20631   }; //i=111 n=1024 twiddle= 7.768885e-01    + i -6.296382e-01
		10'd112: twiddle = { 16'd25329   , -16'd20787   }; //i=112 n=1024 twiddle= 7.730105e-01    + i -6.343933e-01
		10'd113: twiddle = { 16'd25201   , -16'd20942   }; //i=113 n=1024 twiddle= 7.691033e-01    + i -6.391244e-01
		10'd114: twiddle = { 16'd25072   , -16'd21096   }; //i=114 n=1024 twiddle= 7.651673e-01    + i -6.438315e-01
		10'd115: twiddle = { 16'd24942   , -16'd21250   }; //i=115 n=1024 twiddle= 7.612024e-01    + i -6.485144e-01
		10'd116: twiddle = { 16'd24811   , -16'd21403   }; //i=116 n=1024 twiddle= 7.572088e-01    + i -6.531728e-01
		10'd117: twiddle = { 16'd24680   , -16'd21554   }; //i=117 n=1024 twiddle= 7.531868e-01    + i -6.578067e-01
		10'd118: twiddle = { 16'd24547   , -16'd21705   }; //i=118 n=1024 twiddle= 7.491364e-01    + i -6.624158e-01
		10'd119: twiddle = { 16'd24413   , -16'd21856   }; //i=119 n=1024 twiddle= 7.450578e-01    + i -6.669999e-01
		10'd120: twiddle = { 16'd24279   , -16'd22005   }; //i=120 n=1024 twiddle= 7.409511e-01    + i -6.715590e-01
		10'd121: twiddle = { 16'd24143   , -16'd22154   }; //i=121 n=1024 twiddle= 7.368166e-01    + i -6.760927e-01
		10'd122: twiddle = { 16'd24007   , -16'd22301   }; //i=122 n=1024 twiddle= 7.326543e-01    + i -6.806010e-01
		10'd123: twiddle = { 16'd23870   , -16'd22448   }; //i=123 n=1024 twiddle= 7.284644e-01    + i -6.850837e-01
		10'd124: twiddle = { 16'd23731   , -16'd22594   }; //i=124 n=1024 twiddle= 7.242471e-01    + i -6.895405e-01
		10'd125: twiddle = { 16'd23592   , -16'd22739   }; //i=125 n=1024 twiddle= 7.200025e-01    + i -6.939715e-01
		10'd126: twiddle = { 16'd23452   , -16'd22884   }; //i=126 n=1024 twiddle= 7.157308e-01    + i -6.983762e-01
		10'd127: twiddle = { 16'd23311   , -16'd23027   }; //i=127 n=1024 twiddle= 7.114322e-01    + i -7.027547e-01
		10'd128: twiddle = { 16'd23170   , -16'd23170   }; //i=128 n=1024 twiddle= 7.071068e-01    + i -7.071068e-01
		10'd129: twiddle = { 16'd23027   , -16'd23311   }; //i=129 n=1024 twiddle= 7.027547e-01    + i -7.114322e-01
		10'd130: twiddle = { 16'd22884   , -16'd23452   }; //i=130 n=1024 twiddle= 6.983762e-01    + i -7.157308e-01
		10'd131: twiddle = { 16'd22739   , -16'd23592   }; //i=131 n=1024 twiddle= 6.939715e-01    + i -7.200025e-01
		10'd132: twiddle = { 16'd22594   , -16'd23731   }; //i=132 n=1024 twiddle= 6.895405e-01    + i -7.242471e-01
		10'd133: twiddle = { 16'd22448   , -16'd23870   }; //i=133 n=1024 twiddle= 6.850837e-01    + i -7.284644e-01
		10'd134: twiddle = { 16'd22301   , -16'd24007   }; //i=134 n=1024 twiddle= 6.806010e-01    + i -7.326543e-01
		10'd135: twiddle = { 16'd22154   , -16'd24143   }; //i=135 n=1024 twiddle= 6.760927e-01    + i -7.368166e-01
		10'd136: twiddle = { 16'd22005   , -16'd24279   }; //i=136 n=1024 twiddle= 6.715590e-01    + i -7.409511e-01
		10'd137: twiddle = { 16'd21856   , -16'd24413   }; //i=137 n=1024 twiddle= 6.669999e-01    + i -7.450578e-01
		10'd138: twiddle = { 16'd21705   , -16'd24547   }; //i=138 n=1024 twiddle= 6.624158e-01    + i -7.491364e-01
		10'd139: twiddle = { 16'd21554   , -16'd24680   }; //i=139 n=1024 twiddle= 6.578067e-01    + i -7.531868e-01
		10'd140: twiddle = { 16'd21403   , -16'd24811   }; //i=140 n=1024 twiddle= 6.531728e-01    + i -7.572088e-01
		10'd141: twiddle = { 16'd21250   , -16'd24942   }; //i=141 n=1024 twiddle= 6.485144e-01    + i -7.612024e-01
		10'd142: twiddle = { 16'd21096   , -16'd25072   }; //i=142 n=1024 twiddle= 6.438315e-01    + i -7.651673e-01
		10'd143: twiddle = { 16'd20942   , -16'd25201   }; //i=143 n=1024 twiddle= 6.391244e-01    + i -7.691033e-01
		10'd144: twiddle = { 16'd20787   , -16'd25329   }; //i=144 n=1024 twiddle= 6.343933e-01    + i -7.730105e-01
		10'd145: twiddle = { 16'd20631   , -16'd25456   }; //i=145 n=1024 twiddle= 6.296382e-01    + i -7.768885e-01
		10'd146: twiddle = { 16'd20475   , -16'd25582   }; //i=146 n=1024 twiddle= 6.248595e-01    + i -7.807372e-01
		10'd147: twiddle = { 16'd20317   , -16'd25708   }; //i=147 n=1024 twiddle= 6.200572e-01    + i -7.845566e-01
		10'd148: twiddle = { 16'd20159   , -16'd25832   }; //i=148 n=1024 twiddle= 6.152316e-01    + i -7.883464e-01
		10'd149: twiddle = { 16'd20000   , -16'd25955   }; //i=149 n=1024 twiddle= 6.103828e-01    + i -7.921066e-01
		10'd150: twiddle = { 16'd19841   , -16'd26077   }; //i=150 n=1024 twiddle= 6.055110e-01    + i -7.958369e-01
		10'd151: twiddle = { 16'd19680   , -16'd26198   }; //i=151 n=1024 twiddle= 6.006165e-01    + i -7.995373e-01
		10'd152: twiddle = { 16'd19519   , -16'd26319   }; //i=152 n=1024 twiddle= 5.956993e-01    + i -8.032075e-01
		10'd153: twiddle = { 16'd19357   , -16'd26438   }; //i=153 n=1024 twiddle= 5.907597e-01    + i -8.068476e-01
		10'd154: twiddle = { 16'd19195   , -16'd26556   }; //i=154 n=1024 twiddle= 5.857979e-01    + i -8.104572e-01
		10'd155: twiddle = { 16'd19032   , -16'd26674   }; //i=155 n=1024 twiddle= 5.808140e-01    + i -8.140363e-01
		10'd156: twiddle = { 16'd18868   , -16'd26790   }; //i=156 n=1024 twiddle= 5.758082e-01    + i -8.175848e-01
		10'd157: twiddle = { 16'd18703   , -16'd26905   }; //i=157 n=1024 twiddle= 5.707807e-01    + i -8.211025e-01
		10'd158: twiddle = { 16'd18537   , -16'd27019   }; //i=158 n=1024 twiddle= 5.657318e-01    + i -8.245893e-01
		10'd159: twiddle = { 16'd18371   , -16'd27133   }; //i=159 n=1024 twiddle= 5.606616e-01    + i -8.280450e-01
		10'd160: twiddle = { 16'd18204   , -16'd27245   }; //i=160 n=1024 twiddle= 5.555702e-01    + i -8.314696e-01
		10'd161: twiddle = { 16'd18037   , -16'd27356   }; //i=161 n=1024 twiddle= 5.504580e-01    + i -8.348629e-01
		10'd162: twiddle = { 16'd17869   , -16'd27466   }; //i=162 n=1024 twiddle= 5.453250e-01    + i -8.382247e-01
		10'd163: twiddle = { 16'd17700   , -16'd27575   }; //i=163 n=1024 twiddle= 5.401715e-01    + i -8.415550e-01
		10'd164: twiddle = { 16'd17530   , -16'd27683   }; //i=164 n=1024 twiddle= 5.349976e-01    + i -8.448536e-01
		10'd165: twiddle = { 16'd17360   , -16'd27790   }; //i=165 n=1024 twiddle= 5.298036e-01    + i -8.481203e-01
		10'd166: twiddle = { 16'd17189   , -16'd27896   }; //i=166 n=1024 twiddle= 5.245897e-01    + i -8.513552e-01
		10'd167: twiddle = { 16'd17018   , -16'd28001   }; //i=167 n=1024 twiddle= 5.193560e-01    + i -8.545580e-01
		10'd168: twiddle = { 16'd16846   , -16'd28105   }; //i=168 n=1024 twiddle= 5.141027e-01    + i -8.577286e-01
		10'd169: twiddle = { 16'd16673   , -16'd28208   }; //i=169 n=1024 twiddle= 5.088301e-01    + i -8.608669e-01
		10'd170: twiddle = { 16'd16499   , -16'd28310   }; //i=170 n=1024 twiddle= 5.035384e-01    + i -8.639729e-01
		10'd171: twiddle = { 16'd16325   , -16'd28411   }; //i=171 n=1024 twiddle= 4.982277e-01    + i -8.670462e-01
		10'd172: twiddle = { 16'd16151   , -16'd28510   }; //i=172 n=1024 twiddle= 4.928982e-01    + i -8.700870e-01
		10'd173: twiddle = { 16'd15976   , -16'd28609   }; //i=173 n=1024 twiddle= 4.875502e-01    + i -8.730950e-01
		10'd174: twiddle = { 16'd15800   , -16'd28706   }; //i=174 n=1024 twiddle= 4.821838e-01    + i -8.760701e-01
		10'd175: twiddle = { 16'd15623   , -16'd28803   }; //i=175 n=1024 twiddle= 4.767992e-01    + i -8.790122e-01
		10'd176: twiddle = { 16'd15446   , -16'd28898   }; //i=176 n=1024 twiddle= 4.713967e-01    + i -8.819213e-01
		10'd177: twiddle = { 16'd15269   , -16'd28992   }; //i=177 n=1024 twiddle= 4.659765e-01    + i -8.847971e-01
		10'd178: twiddle = { 16'd15090   , -16'd29085   }; //i=178 n=1024 twiddle= 4.605387e-01    + i -8.876396e-01
		10'd179: twiddle = { 16'd14912   , -16'd29177   }; //i=179 n=1024 twiddle= 4.550836e-01    + i -8.904487e-01
		10'd180: twiddle = { 16'd14732   , -16'd29268   }; //i=180 n=1024 twiddle= 4.496113e-01    + i -8.932243e-01
		10'd181: twiddle = { 16'd14553   , -16'd29358   }; //i=181 n=1024 twiddle= 4.441221e-01    + i -8.959662e-01
		10'd182: twiddle = { 16'd14372   , -16'd29447   }; //i=182 n=1024 twiddle= 4.386162e-01    + i -8.986745e-01
		10'd183: twiddle = { 16'd14191   , -16'd29534   }; //i=183 n=1024 twiddle= 4.330938e-01    + i -9.013488e-01
		10'd184: twiddle = { 16'd14010   , -16'd29621   }; //i=184 n=1024 twiddle= 4.275551e-01    + i -9.039893e-01
		10'd185: twiddle = { 16'd13828   , -16'd29706   }; //i=185 n=1024 twiddle= 4.220003e-01    + i -9.065957e-01
		10'd186: twiddle = { 16'd13645   , -16'd29791   }; //i=186 n=1024 twiddle= 4.164296e-01    + i -9.091680e-01
		10'd187: twiddle = { 16'd13462   , -16'd29874   }; //i=187 n=1024 twiddle= 4.108432e-01    + i -9.117060e-01
		10'd188: twiddle = { 16'd13279   , -16'd29956   }; //i=188 n=1024 twiddle= 4.052413e-01    + i -9.142098e-01
		10'd189: twiddle = { 16'd13094   , -16'd30037   }; //i=189 n=1024 twiddle= 3.996242e-01    + i -9.166791e-01
		10'd190: twiddle = { 16'd12910   , -16'd30117   }; //i=190 n=1024 twiddle= 3.939920e-01    + i -9.191139e-01
		10'd191: twiddle = { 16'd12725   , -16'd30195   }; //i=191 n=1024 twiddle= 3.883450e-01    + i -9.215140e-01
		10'd192: twiddle = { 16'd12539   , -16'd30273   }; //i=192 n=1024 twiddle= 3.826834e-01    + i -9.238795e-01
		10'd193: twiddle = { 16'd12353   , -16'd30349   }; //i=193 n=1024 twiddle= 3.770074e-01    + i -9.262102e-01
		10'd194: twiddle = { 16'd12167   , -16'd30424   }; //i=194 n=1024 twiddle= 3.713172e-01    + i -9.285061e-01
		10'd195: twiddle = { 16'd11980   , -16'd30498   }; //i=195 n=1024 twiddle= 3.656130e-01    + i -9.307670e-01
		10'd196: twiddle = { 16'd11793   , -16'd30571   }; //i=196 n=1024 twiddle= 3.598950e-01    + i -9.329928e-01
		10'd197: twiddle = { 16'd11605   , -16'd30643   }; //i=197 n=1024 twiddle= 3.541635e-01    + i -9.351835e-01
		10'd198: twiddle = { 16'd11417   , -16'd30714   }; //i=198 n=1024 twiddle= 3.484187e-01    + i -9.373390e-01
		10'd199: twiddle = { 16'd11228   , -16'd30783   }; //i=199 n=1024 twiddle= 3.426607e-01    + i -9.394592e-01
		10'd200: twiddle = { 16'd11039   , -16'd30852   }; //i=200 n=1024 twiddle= 3.368899e-01    + i -9.415441e-01
		10'd201: twiddle = { 16'd10849   , -16'd30919   }; //i=201 n=1024 twiddle= 3.311063e-01    + i -9.435935e-01
		10'd202: twiddle = { 16'd10659   , -16'd30985   }; //i=202 n=1024 twiddle= 3.253103e-01    + i -9.456073e-01
		10'd203: twiddle = { 16'd10469   , -16'd31050   }; //i=203 n=1024 twiddle= 3.195020e-01    + i -9.475856e-01
		10'd204: twiddle = { 16'd10278   , -16'd31113   }; //i=204 n=1024 twiddle= 3.136817e-01    + i -9.495282e-01
		10'd205: twiddle = { 16'd10087   , -16'd31176   }; //i=205 n=1024 twiddle= 3.078496e-01    + i -9.514350e-01
		10'd206: twiddle = { 16'd9896    , -16'd31237   }; //i=206 n=1024 twiddle= 3.020059e-01    + i -9.533060e-01
		10'd207: twiddle = { 16'd9704    , -16'd31297   }; //i=207 n=1024 twiddle= 2.961509e-01    + i -9.551412e-01
		10'd208: twiddle = { 16'd9512    , -16'd31356   }; //i=208 n=1024 twiddle= 2.902847e-01    + i -9.569403e-01
		10'd209: twiddle = { 16'd9319    , -16'd31414   }; //i=209 n=1024 twiddle= 2.844075e-01    + i -9.587035e-01
		10'd210: twiddle = { 16'd9126    , -16'd31470   }; //i=210 n=1024 twiddle= 2.785197e-01    + i -9.604305e-01
		10'd211: twiddle = { 16'd8933    , -16'd31526   }; //i=211 n=1024 twiddle= 2.726214e-01    + i -9.621214e-01
		10'd212: twiddle = { 16'd8739    , -16'd31580   }; //i=212 n=1024 twiddle= 2.667128e-01    + i -9.637761e-01
		10'd213: twiddle = { 16'd8545    , -16'd31633   }; //i=213 n=1024 twiddle= 2.607941e-01    + i -9.653944e-01
		10'd214: twiddle = { 16'd8351    , -16'd31685   }; //i=214 n=1024 twiddle= 2.548657e-01    + i -9.669765e-01
		10'd215: twiddle = { 16'd8157    , -16'd31736   }; //i=215 n=1024 twiddle= 2.489276e-01    + i -9.685221e-01
		10'd216: twiddle = { 16'd7962    , -16'd31785   }; //i=216 n=1024 twiddle= 2.429802e-01    + i -9.700313e-01
		10'd217: twiddle = { 16'd7767    , -16'd31833   }; //i=217 n=1024 twiddle= 2.370236e-01    + i -9.715039e-01
		10'd218: twiddle = { 16'd7571    , -16'd31880   }; //i=218 n=1024 twiddle= 2.310581e-01    + i -9.729400e-01
		10'd219: twiddle = { 16'd7375    , -16'd31926   }; //i=219 n=1024 twiddle= 2.250839e-01    + i -9.743394e-01
		10'd220: twiddle = { 16'd7179    , -16'd31971   }; //i=220 n=1024 twiddle= 2.191012e-01    + i -9.757021e-01
		10'd221: twiddle = { 16'd6983    , -16'd32014   }; //i=221 n=1024 twiddle= 2.131103e-01    + i -9.770281e-01
		10'd222: twiddle = { 16'd6786    , -16'd32057   }; //i=222 n=1024 twiddle= 2.071114e-01    + i -9.783174e-01
		10'd223: twiddle = { 16'd6590    , -16'd32098   }; //i=223 n=1024 twiddle= 2.011046e-01    + i -9.795698e-01
		10'd224: twiddle = { 16'd6393    , -16'd32137   }; //i=224 n=1024 twiddle= 1.950903e-01    + i -9.807853e-01
		10'd225: twiddle = { 16'd6195    , -16'd32176   }; //i=225 n=1024 twiddle= 1.890687e-01    + i -9.819639e-01
		10'd226: twiddle = { 16'd5998    , -16'd32213   }; //i=226 n=1024 twiddle= 1.830399e-01    + i -9.831055e-01
		10'd227: twiddle = { 16'd5800    , -16'd32250   }; //i=227 n=1024 twiddle= 1.770042e-01    + i -9.842101e-01
		10'd228: twiddle = { 16'd5602    , -16'd32285   }; //i=228 n=1024 twiddle= 1.709619e-01    + i -9.852776e-01
		10'd229: twiddle = { 16'd5404    , -16'd32318   }; //i=229 n=1024 twiddle= 1.649131e-01    + i -9.863081e-01
		10'd230: twiddle = { 16'd5205    , -16'd32351   }; //i=230 n=1024 twiddle= 1.588581e-01    + i -9.873014e-01
		10'd231: twiddle = { 16'd5007    , -16'd32382   }; //i=231 n=1024 twiddle= 1.527972e-01    + i -9.882576e-01
		10'd232: twiddle = { 16'd4808    , -16'd32412   }; //i=232 n=1024 twiddle= 1.467305e-01    + i -9.891765e-01
		10'd233: twiddle = { 16'd4609    , -16'd32441   }; //i=233 n=1024 twiddle= 1.406582e-01    + i -9.900582e-01
		10'd234: twiddle = { 16'd4410    , -16'd32469   }; //i=234 n=1024 twiddle= 1.345807e-01    + i -9.909026e-01
		10'd235: twiddle = { 16'd4210    , -16'd32495   }; //i=235 n=1024 twiddle= 1.284981e-01    + i -9.917098e-01
		10'd236: twiddle = { 16'd4011    , -16'd32521   }; //i=236 n=1024 twiddle= 1.224107e-01    + i -9.924795e-01
		10'd237: twiddle = { 16'd3811    , -16'd32545   }; //i=237 n=1024 twiddle= 1.163186e-01    + i -9.932119e-01
		10'd238: twiddle = { 16'd3612    , -16'd32567   }; //i=238 n=1024 twiddle= 1.102222e-01    + i -9.939070e-01
		10'd239: twiddle = { 16'd3412    , -16'd32589   }; //i=239 n=1024 twiddle= 1.041216e-01    + i -9.945646e-01
		10'd240: twiddle = { 16'd3212    , -16'd32609   }; //i=240 n=1024 twiddle= 9.801714e-02    + i -9.951847e-01
		10'd241: twiddle = { 16'd3012    , -16'd32628   }; //i=241 n=1024 twiddle= 9.190896e-02    + i -9.957674e-01
		10'd242: twiddle = { 16'd2811    , -16'd32646   }; //i=242 n=1024 twiddle= 8.579731e-02    + i -9.963126e-01
		10'd243: twiddle = { 16'd2611    , -16'd32663   }; //i=243 n=1024 twiddle= 7.968244e-02    + i -9.968203e-01
		10'd244: twiddle = { 16'd2410    , -16'd32678   }; //i=244 n=1024 twiddle= 7.356456e-02    + i -9.972905e-01
		10'd245: twiddle = { 16'd2210    , -16'd32692   }; //i=245 n=1024 twiddle= 6.744392e-02    + i -9.977231e-01
		10'd246: twiddle = { 16'd2009    , -16'd32705   }; //i=246 n=1024 twiddle= 6.132074e-02    + i -9.981181e-01
		10'd247: twiddle = { 16'd1809    , -16'd32717   }; //i=247 n=1024 twiddle= 5.519524e-02    + i -9.984756e-01
		10'd248: twiddle = { 16'd1608    , -16'd32728   }; //i=248 n=1024 twiddle= 4.906767e-02    + i -9.987955e-01
		10'd249: twiddle = { 16'd1407    , -16'd32737   }; //i=249 n=1024 twiddle= 4.293826e-02    + i -9.990777e-01
		10'd250: twiddle = { 16'd1206    , -16'd32745   }; //i=250 n=1024 twiddle= 3.680722e-02    + i -9.993224e-01
		10'd251: twiddle = { 16'd1005    , -16'd32752   }; //i=251 n=1024 twiddle= 3.067480e-02    + i -9.995294e-01
		10'd252: twiddle = { 16'd804     , -16'd32757   }; //i=252 n=1024 twiddle= 2.454123e-02    + i -9.996988e-01
		10'd253: twiddle = { 16'd603     , -16'd32761   }; //i=253 n=1024 twiddle= 1.840673e-02    + i -9.998306e-01
		10'd254: twiddle = { 16'd402     , -16'd32765   }; //i=254 n=1024 twiddle= 1.227154e-02    + i -9.999247e-01
		10'd255: twiddle = { 16'd201     , -16'd32766   }; //i=255 n=1024 twiddle= 6.135885e-03    + i -9.999812e-01
		10'd256: twiddle = { 16'd0       , -16'd32767   }; //i=256 n=1024 twiddle= 6.123234e-17    + i -1
		10'd257: twiddle = {-16'd201     , -16'd32766   }; //i=257 n=1024 twiddle= -6.135885e-03   + i -9.999812e-01
		10'd258: twiddle = {-16'd402     , -16'd32765   }; //i=258 n=1024 twiddle= -1.227154e-02   + i -9.999247e-01
		10'd259: twiddle = {-16'd603     , -16'd32761   }; //i=259 n=1024 twiddle= -1.840673e-02   + i -9.998306e-01
		10'd260: twiddle = {-16'd804     , -16'd32757   }; //i=260 n=1024 twiddle= -2.454123e-02   + i -9.996988e-01
		10'd261: twiddle = {-16'd1005    , -16'd32752   }; //i=261 n=1024 twiddle= -3.067480e-02   + i -9.995294e-01
		10'd262: twiddle = {-16'd1206    , -16'd32745   }; //i=262 n=1024 twiddle= -3.680722e-02   + i -9.993224e-01
		10'd263: twiddle = {-16'd1407    , -16'd32737   }; //i=263 n=1024 twiddle= -4.293826e-02   + i -9.990777e-01
		10'd264: twiddle = {-16'd1608    , -16'd32728   }; //i=264 n=1024 twiddle= -4.906767e-02   + i -9.987955e-01
		10'd265: twiddle = {-16'd1809    , -16'd32717   }; //i=265 n=1024 twiddle= -5.519524e-02   + i -9.984756e-01
		10'd266: twiddle = {-16'd2009    , -16'd32705   }; //i=266 n=1024 twiddle= -6.132074e-02   + i -9.981181e-01
		10'd267: twiddle = {-16'd2210    , -16'd32692   }; //i=267 n=1024 twiddle= -6.744392e-02   + i -9.977231e-01
		10'd268: twiddle = {-16'd2410    , -16'd32678   }; //i=268 n=1024 twiddle= -7.356456e-02   + i -9.972905e-01
		10'd269: twiddle = {-16'd2611    , -16'd32663   }; //i=269 n=1024 twiddle= -7.968244e-02   + i -9.968203e-01
		10'd270: twiddle = {-16'd2811    , -16'd32646   }; //i=270 n=1024 twiddle= -8.579731e-02   + i -9.963126e-01
		10'd271: twiddle = {-16'd3012    , -16'd32628   }; //i=271 n=1024 twiddle= -9.190896e-02   + i -9.957674e-01
		10'd272: twiddle = {-16'd3212    , -16'd32609   }; //i=272 n=1024 twiddle= -9.801714e-02   + i -9.951847e-01
		10'd273: twiddle = {-16'd3412    , -16'd32589   }; //i=273 n=1024 twiddle= -1.041216e-01   + i -9.945646e-01
		10'd274: twiddle = {-16'd3612    , -16'd32567   }; //i=274 n=1024 twiddle= -1.102222e-01   + i -9.939070e-01
		10'd275: twiddle = {-16'd3811    , -16'd32545   }; //i=275 n=1024 twiddle= -1.163186e-01   + i -9.932119e-01
		10'd276: twiddle = {-16'd4011    , -16'd32521   }; //i=276 n=1024 twiddle= -1.224107e-01   + i -9.924795e-01
		10'd277: twiddle = {-16'd4210    , -16'd32495   }; //i=277 n=1024 twiddle= -1.284981e-01   + i -9.917098e-01
		10'd278: twiddle = {-16'd4410    , -16'd32469   }; //i=278 n=1024 twiddle= -1.345807e-01   + i -9.909026e-01
		10'd279: twiddle = {-16'd4609    , -16'd32441   }; //i=279 n=1024 twiddle= -1.406582e-01   + i -9.900582e-01
		10'd280: twiddle = {-16'd4808    , -16'd32412   }; //i=280 n=1024 twiddle= -1.467305e-01   + i -9.891765e-01
		10'd281: twiddle = {-16'd5007    , -16'd32382   }; //i=281 n=1024 twiddle= -1.527972e-01   + i -9.882576e-01
		10'd282: twiddle = {-16'd5205    , -16'd32351   }; //i=282 n=1024 twiddle= -1.588581e-01   + i -9.873014e-01
		10'd283: twiddle = {-16'd5404    , -16'd32318   }; //i=283 n=1024 twiddle= -1.649131e-01   + i -9.863081e-01
		10'd284: twiddle = {-16'd5602    , -16'd32285   }; //i=284 n=1024 twiddle= -1.709619e-01   + i -9.852776e-01
		10'd285: twiddle = {-16'd5800    , -16'd32250   }; //i=285 n=1024 twiddle= -1.770042e-01   + i -9.842101e-01
		10'd286: twiddle = {-16'd5998    , -16'd32213   }; //i=286 n=1024 twiddle= -1.830399e-01   + i -9.831055e-01
		10'd287: twiddle = {-16'd6195    , -16'd32176   }; //i=287 n=1024 twiddle= -1.890687e-01   + i -9.819639e-01
		10'd288: twiddle = {-16'd6393    , -16'd32137   }; //i=288 n=1024 twiddle= -1.950903e-01   + i -9.807853e-01
		10'd289: twiddle = {-16'd6590    , -16'd32098   }; //i=289 n=1024 twiddle= -2.011046e-01   + i -9.795698e-01
		10'd290: twiddle = {-16'd6786    , -16'd32057   }; //i=290 n=1024 twiddle= -2.071114e-01   + i -9.783174e-01
		10'd291: twiddle = {-16'd6983    , -16'd32014   }; //i=291 n=1024 twiddle= -2.131103e-01   + i -9.770281e-01
		10'd292: twiddle = {-16'd7179    , -16'd31971   }; //i=292 n=1024 twiddle= -2.191012e-01   + i -9.757021e-01
		10'd293: twiddle = {-16'd7375    , -16'd31926   }; //i=293 n=1024 twiddle= -2.250839e-01   + i -9.743394e-01
		10'd294: twiddle = {-16'd7571    , -16'd31880   }; //i=294 n=1024 twiddle= -2.310581e-01   + i -9.729400e-01
		10'd295: twiddle = {-16'd7767    , -16'd31833   }; //i=295 n=1024 twiddle= -2.370236e-01   + i -9.715039e-01
		10'd296: twiddle = {-16'd7962    , -16'd31785   }; //i=296 n=1024 twiddle= -2.429802e-01   + i -9.700313e-01
		10'd297: twiddle = {-16'd8157    , -16'd31736   }; //i=297 n=1024 twiddle= -2.489276e-01   + i -9.685221e-01
		10'd298: twiddle = {-16'd8351    , -16'd31685   }; //i=298 n=1024 twiddle= -2.548657e-01   + i -9.669765e-01
		10'd299: twiddle = {-16'd8545    , -16'd31633   }; //i=299 n=1024 twiddle= -2.607941e-01   + i -9.653944e-01
		10'd300: twiddle = {-16'd8739    , -16'd31580   }; //i=300 n=1024 twiddle= -2.667128e-01   + i -9.637761e-01
		10'd301: twiddle = {-16'd8933    , -16'd31526   }; //i=301 n=1024 twiddle= -2.726214e-01   + i -9.621214e-01
		10'd302: twiddle = {-16'd9126    , -16'd31470   }; //i=302 n=1024 twiddle= -2.785197e-01   + i -9.604305e-01
		10'd303: twiddle = {-16'd9319    , -16'd31414   }; //i=303 n=1024 twiddle= -2.844075e-01   + i -9.587035e-01
		10'd304: twiddle = {-16'd9512    , -16'd31356   }; //i=304 n=1024 twiddle= -2.902847e-01   + i -9.569403e-01
		10'd305: twiddle = {-16'd9704    , -16'd31297   }; //i=305 n=1024 twiddle= -2.961509e-01   + i -9.551412e-01
		10'd306: twiddle = {-16'd9896    , -16'd31237   }; //i=306 n=1024 twiddle= -3.020059e-01   + i -9.533060e-01
		10'd307: twiddle = {-16'd10087   , -16'd31176   }; //i=307 n=1024 twiddle= -3.078496e-01   + i -9.514350e-01
		10'd308: twiddle = {-16'd10278   , -16'd31113   }; //i=308 n=1024 twiddle= -3.136817e-01   + i -9.495282e-01
		10'd309: twiddle = {-16'd10469   , -16'd31050   }; //i=309 n=1024 twiddle= -3.195020e-01   + i -9.475856e-01
		10'd310: twiddle = {-16'd10659   , -16'd30985   }; //i=310 n=1024 twiddle= -3.253103e-01   + i -9.456073e-01
		10'd311: twiddle = {-16'd10849   , -16'd30919   }; //i=311 n=1024 twiddle= -3.311063e-01   + i -9.435935e-01
		10'd312: twiddle = {-16'd11039   , -16'd30852   }; //i=312 n=1024 twiddle= -3.368899e-01   + i -9.415441e-01
		10'd313: twiddle = {-16'd11228   , -16'd30783   }; //i=313 n=1024 twiddle= -3.426607e-01   + i -9.394592e-01
		10'd314: twiddle = {-16'd11417   , -16'd30714   }; //i=314 n=1024 twiddle= -3.484187e-01   + i -9.373390e-01
		10'd315: twiddle = {-16'd11605   , -16'd30643   }; //i=315 n=1024 twiddle= -3.541635e-01   + i -9.351835e-01
		10'd316: twiddle = {-16'd11793   , -16'd30571   }; //i=316 n=1024 twiddle= -3.598950e-01   + i -9.329928e-01
		10'd317: twiddle = {-16'd11980   , -16'd30498   }; //i=317 n=1024 twiddle= -3.656130e-01   + i -9.307670e-01
		10'd318: twiddle = {-16'd12167   , -16'd30424   }; //i=318 n=1024 twiddle= -3.713172e-01   + i -9.285061e-01
		10'd319: twiddle = {-16'd12353   , -16'd30349   }; //i=319 n=1024 twiddle= -3.770074e-01   + i -9.262102e-01
		10'd320: twiddle = {-16'd12539   , -16'd30273   }; //i=320 n=1024 twiddle= -3.826834e-01   + i -9.238795e-01
		10'd321: twiddle = {-16'd12725   , -16'd30195   }; //i=321 n=1024 twiddle= -3.883450e-01   + i -9.215140e-01
		10'd322: twiddle = {-16'd12910   , -16'd30117   }; //i=322 n=1024 twiddle= -3.939920e-01   + i -9.191139e-01
		10'd323: twiddle = {-16'd13094   , -16'd30037   }; //i=323 n=1024 twiddle= -3.996242e-01   + i -9.166791e-01
		10'd324: twiddle = {-16'd13279   , -16'd29956   }; //i=324 n=1024 twiddle= -4.052413e-01   + i -9.142098e-01
		10'd325: twiddle = {-16'd13462   , -16'd29874   }; //i=325 n=1024 twiddle= -4.108432e-01   + i -9.117060e-01
		10'd326: twiddle = {-16'd13645   , -16'd29791   }; //i=326 n=1024 twiddle= -4.164296e-01   + i -9.091680e-01
		10'd327: twiddle = {-16'd13828   , -16'd29706   }; //i=327 n=1024 twiddle= -4.220003e-01   + i -9.065957e-01
		10'd328: twiddle = {-16'd14010   , -16'd29621   }; //i=328 n=1024 twiddle= -4.275551e-01   + i -9.039893e-01
		10'd329: twiddle = {-16'd14191   , -16'd29534   }; //i=329 n=1024 twiddle= -4.330938e-01   + i -9.013488e-01
		10'd330: twiddle = {-16'd14372   , -16'd29447   }; //i=330 n=1024 twiddle= -4.386162e-01   + i -8.986745e-01
		10'd331: twiddle = {-16'd14553   , -16'd29358   }; //i=331 n=1024 twiddle= -4.441221e-01   + i -8.959662e-01
		10'd332: twiddle = {-16'd14732   , -16'd29268   }; //i=332 n=1024 twiddle= -4.496113e-01   + i -8.932243e-01
		10'd333: twiddle = {-16'd14912   , -16'd29177   }; //i=333 n=1024 twiddle= -4.550836e-01   + i -8.904487e-01
		10'd334: twiddle = {-16'd15090   , -16'd29085   }; //i=334 n=1024 twiddle= -4.605387e-01   + i -8.876396e-01
		10'd335: twiddle = {-16'd15269   , -16'd28992   }; //i=335 n=1024 twiddle= -4.659765e-01   + i -8.847971e-01
		10'd336: twiddle = {-16'd15446   , -16'd28898   }; //i=336 n=1024 twiddle= -4.713967e-01   + i -8.819213e-01
		10'd337: twiddle = {-16'd15623   , -16'd28803   }; //i=337 n=1024 twiddle= -4.767992e-01   + i -8.790122e-01
		10'd338: twiddle = {-16'd15800   , -16'd28706   }; //i=338 n=1024 twiddle= -4.821838e-01   + i -8.760701e-01
		10'd339: twiddle = {-16'd15976   , -16'd28609   }; //i=339 n=1024 twiddle= -4.875502e-01   + i -8.730950e-01
		10'd340: twiddle = {-16'd16151   , -16'd28510   }; //i=340 n=1024 twiddle= -4.928982e-01   + i -8.700870e-01
		10'd341: twiddle = {-16'd16325   , -16'd28411   }; //i=341 n=1024 twiddle= -4.982277e-01   + i -8.670462e-01
		10'd342: twiddle = {-16'd16499   , -16'd28310   }; //i=342 n=1024 twiddle= -5.035384e-01   + i -8.639729e-01
		10'd343: twiddle = {-16'd16673   , -16'd28208   }; //i=343 n=1024 twiddle= -5.088301e-01   + i -8.608669e-01
		10'd344: twiddle = {-16'd16846   , -16'd28105   }; //i=344 n=1024 twiddle= -5.141027e-01   + i -8.577286e-01
		10'd345: twiddle = {-16'd17018   , -16'd28001   }; //i=345 n=1024 twiddle= -5.193560e-01   + i -8.545580e-01
		10'd346: twiddle = {-16'd17189   , -16'd27896   }; //i=346 n=1024 twiddle= -5.245897e-01   + i -8.513552e-01
		10'd347: twiddle = {-16'd17360   , -16'd27790   }; //i=347 n=1024 twiddle= -5.298036e-01   + i -8.481203e-01
		10'd348: twiddle = {-16'd17530   , -16'd27683   }; //i=348 n=1024 twiddle= -5.349976e-01   + i -8.448536e-01
		10'd349: twiddle = {-16'd17700   , -16'd27575   }; //i=349 n=1024 twiddle= -5.401715e-01   + i -8.415550e-01
		10'd350: twiddle = {-16'd17869   , -16'd27466   }; //i=350 n=1024 twiddle= -5.453250e-01   + i -8.382247e-01
		10'd351: twiddle = {-16'd18037   , -16'd27356   }; //i=351 n=1024 twiddle= -5.504580e-01   + i -8.348629e-01
		10'd352: twiddle = {-16'd18204   , -16'd27245   }; //i=352 n=1024 twiddle= -5.555702e-01   + i -8.314696e-01
		10'd353: twiddle = {-16'd18371   , -16'd27133   }; //i=353 n=1024 twiddle= -5.606616e-01   + i -8.280450e-01
		10'd354: twiddle = {-16'd18537   , -16'd27019   }; //i=354 n=1024 twiddle= -5.657318e-01   + i -8.245893e-01
		10'd355: twiddle = {-16'd18703   , -16'd26905   }; //i=355 n=1024 twiddle= -5.707807e-01   + i -8.211025e-01
		10'd356: twiddle = {-16'd18868   , -16'd26790   }; //i=356 n=1024 twiddle= -5.758082e-01   + i -8.175848e-01
		10'd357: twiddle = {-16'd19032   , -16'd26674   }; //i=357 n=1024 twiddle= -5.808140e-01   + i -8.140363e-01
		10'd358: twiddle = {-16'd19195   , -16'd26556   }; //i=358 n=1024 twiddle= -5.857979e-01   + i -8.104572e-01
		10'd359: twiddle = {-16'd19357   , -16'd26438   }; //i=359 n=1024 twiddle= -5.907597e-01   + i -8.068476e-01
		10'd360: twiddle = {-16'd19519   , -16'd26319   }; //i=360 n=1024 twiddle= -5.956993e-01   + i -8.032075e-01
		10'd361: twiddle = {-16'd19680   , -16'd26198   }; //i=361 n=1024 twiddle= -6.006165e-01   + i -7.995373e-01
		10'd362: twiddle = {-16'd19841   , -16'd26077   }; //i=362 n=1024 twiddle= -6.055110e-01   + i -7.958369e-01
		10'd363: twiddle = {-16'd20000   , -16'd25955   }; //i=363 n=1024 twiddle= -6.103828e-01   + i -7.921066e-01
		10'd364: twiddle = {-16'd20159   , -16'd25832   }; //i=364 n=1024 twiddle= -6.152316e-01   + i -7.883464e-01
		10'd365: twiddle = {-16'd20317   , -16'd25708   }; //i=365 n=1024 twiddle= -6.200572e-01   + i -7.845566e-01
		10'd366: twiddle = {-16'd20475   , -16'd25582   }; //i=366 n=1024 twiddle= -6.248595e-01   + i -7.807372e-01
		10'd367: twiddle = {-16'd20631   , -16'd25456   }; //i=367 n=1024 twiddle= -6.296382e-01   + i -7.768885e-01
		10'd368: twiddle = {-16'd20787   , -16'd25329   }; //i=368 n=1024 twiddle= -6.343933e-01   + i -7.730105e-01
		10'd369: twiddle = {-16'd20942   , -16'd25201   }; //i=369 n=1024 twiddle= -6.391244e-01   + i -7.691033e-01
		10'd370: twiddle = {-16'd21096   , -16'd25072   }; //i=370 n=1024 twiddle= -6.438315e-01   + i -7.651673e-01
		10'd371: twiddle = {-16'd21250   , -16'd24942   }; //i=371 n=1024 twiddle= -6.485144e-01   + i -7.612024e-01
		10'd372: twiddle = {-16'd21403   , -16'd24811   }; //i=372 n=1024 twiddle= -6.531728e-01   + i -7.572088e-01
		10'd373: twiddle = {-16'd21554   , -16'd24680   }; //i=373 n=1024 twiddle= -6.578067e-01   + i -7.531868e-01
		10'd374: twiddle = {-16'd21705   , -16'd24547   }; //i=374 n=1024 twiddle= -6.624158e-01   + i -7.491364e-01
		10'd375: twiddle = {-16'd21856   , -16'd24413   }; //i=375 n=1024 twiddle= -6.669999e-01   + i -7.450578e-01
		10'd376: twiddle = {-16'd22005   , -16'd24279   }; //i=376 n=1024 twiddle= -6.715590e-01   + i -7.409511e-01
		10'd377: twiddle = {-16'd22154   , -16'd24143   }; //i=377 n=1024 twiddle= -6.760927e-01   + i -7.368166e-01
		10'd378: twiddle = {-16'd22301   , -16'd24007   }; //i=378 n=1024 twiddle= -6.806010e-01   + i -7.326543e-01
		10'd379: twiddle = {-16'd22448   , -16'd23870   }; //i=379 n=1024 twiddle= -6.850837e-01   + i -7.284644e-01
		10'd380: twiddle = {-16'd22594   , -16'd23731   }; //i=380 n=1024 twiddle= -6.895405e-01   + i -7.242471e-01
		10'd381: twiddle = {-16'd22739   , -16'd23592   }; //i=381 n=1024 twiddle= -6.939715e-01   + i -7.200025e-01
		10'd382: twiddle = {-16'd22884   , -16'd23452   }; //i=382 n=1024 twiddle= -6.983762e-01   + i -7.157308e-01
		10'd383: twiddle = {-16'd23027   , -16'd23311   }; //i=383 n=1024 twiddle= -7.027547e-01   + i -7.114322e-01
		10'd384: twiddle = {-16'd23170   , -16'd23170   }; //i=384 n=1024 twiddle= -7.071068e-01   + i -7.071068e-01
		10'd385: twiddle = {-16'd23311   , -16'd23027   }; //i=385 n=1024 twiddle= -7.114322e-01   + i -7.027547e-01
		10'd386: twiddle = {-16'd23452   , -16'd22884   }; //i=386 n=1024 twiddle= -7.157308e-01   + i -6.983762e-01
		10'd387: twiddle = {-16'd23592   , -16'd22739   }; //i=387 n=1024 twiddle= -7.200025e-01   + i -6.939715e-01
		10'd388: twiddle = {-16'd23731   , -16'd22594   }; //i=388 n=1024 twiddle= -7.242471e-01   + i -6.895405e-01
		10'd389: twiddle = {-16'd23870   , -16'd22448   }; //i=389 n=1024 twiddle= -7.284644e-01   + i -6.850837e-01
		10'd390: twiddle = {-16'd24007   , -16'd22301   }; //i=390 n=1024 twiddle= -7.326543e-01   + i -6.806010e-01
		10'd391: twiddle = {-16'd24143   , -16'd22154   }; //i=391 n=1024 twiddle= -7.368166e-01   + i -6.760927e-01
		10'd392: twiddle = {-16'd24279   , -16'd22005   }; //i=392 n=1024 twiddle= -7.409511e-01   + i -6.715590e-01
		10'd393: twiddle = {-16'd24413   , -16'd21856   }; //i=393 n=1024 twiddle= -7.450578e-01   + i -6.669999e-01
		10'd394: twiddle = {-16'd24547   , -16'd21705   }; //i=394 n=1024 twiddle= -7.491364e-01   + i -6.624158e-01
		10'd395: twiddle = {-16'd24680   , -16'd21554   }; //i=395 n=1024 twiddle= -7.531868e-01   + i -6.578067e-01
		10'd396: twiddle = {-16'd24811   , -16'd21403   }; //i=396 n=1024 twiddle= -7.572088e-01   + i -6.531728e-01
		10'd397: twiddle = {-16'd24942   , -16'd21250   }; //i=397 n=1024 twiddle= -7.612024e-01   + i -6.485144e-01
		10'd398: twiddle = {-16'd25072   , -16'd21096   }; //i=398 n=1024 twiddle= -7.651673e-01   + i -6.438315e-01
		10'd399: twiddle = {-16'd25201   , -16'd20942   }; //i=399 n=1024 twiddle= -7.691033e-01   + i -6.391244e-01
		10'd400: twiddle = {-16'd25329   , -16'd20787   }; //i=400 n=1024 twiddle= -7.730105e-01   + i -6.343933e-01
		10'd401: twiddle = {-16'd25456   , -16'd20631   }; //i=401 n=1024 twiddle= -7.768885e-01   + i -6.296382e-01
		10'd402: twiddle = {-16'd25582   , -16'd20475   }; //i=402 n=1024 twiddle= -7.807372e-01   + i -6.248595e-01
		10'd403: twiddle = {-16'd25708   , -16'd20317   }; //i=403 n=1024 twiddle= -7.845566e-01   + i -6.200572e-01
		10'd404: twiddle = {-16'd25832   , -16'd20159   }; //i=404 n=1024 twiddle= -7.883464e-01   + i -6.152316e-01
		10'd405: twiddle = {-16'd25955   , -16'd20000   }; //i=405 n=1024 twiddle= -7.921066e-01   + i -6.103828e-01
		10'd406: twiddle = {-16'd26077   , -16'd19841   }; //i=406 n=1024 twiddle= -7.958369e-01   + i -6.055110e-01
		10'd407: twiddle = {-16'd26198   , -16'd19680   }; //i=407 n=1024 twiddle= -7.995373e-01   + i -6.006165e-01
		10'd408: twiddle = {-16'd26319   , -16'd19519   }; //i=408 n=1024 twiddle= -8.032075e-01   + i -5.956993e-01
		10'd409: twiddle = {-16'd26438   , -16'd19357   }; //i=409 n=1024 twiddle= -8.068476e-01   + i -5.907597e-01
		10'd410: twiddle = {-16'd26556   , -16'd19195   }; //i=410 n=1024 twiddle= -8.104572e-01   + i -5.857979e-01
		10'd411: twiddle = {-16'd26674   , -16'd19032   }; //i=411 n=1024 twiddle= -8.140363e-01   + i -5.808140e-01
		10'd412: twiddle = {-16'd26790   , -16'd18868   }; //i=412 n=1024 twiddle= -8.175848e-01   + i -5.758082e-01
		10'd413: twiddle = {-16'd26905   , -16'd18703   }; //i=413 n=1024 twiddle= -8.211025e-01   + i -5.707807e-01
		10'd414: twiddle = {-16'd27019   , -16'd18537   }; //i=414 n=1024 twiddle= -8.245893e-01   + i -5.657318e-01
		10'd415: twiddle = {-16'd27133   , -16'd18371   }; //i=415 n=1024 twiddle= -8.280450e-01   + i -5.606616e-01
		10'd416: twiddle = {-16'd27245   , -16'd18204   }; //i=416 n=1024 twiddle= -8.314696e-01   + i -5.555702e-01
		10'd417: twiddle = {-16'd27356   , -16'd18037   }; //i=417 n=1024 twiddle= -8.348629e-01   + i -5.504580e-01
		10'd418: twiddle = {-16'd27466   , -16'd17869   }; //i=418 n=1024 twiddle= -8.382247e-01   + i -5.453250e-01
		10'd419: twiddle = {-16'd27575   , -16'd17700   }; //i=419 n=1024 twiddle= -8.415550e-01   + i -5.401715e-01
		10'd420: twiddle = {-16'd27683   , -16'd17530   }; //i=420 n=1024 twiddle= -8.448536e-01   + i -5.349976e-01
		10'd421: twiddle = {-16'd27790   , -16'd17360   }; //i=421 n=1024 twiddle= -8.481203e-01   + i -5.298036e-01
		10'd422: twiddle = {-16'd27896   , -16'd17189   }; //i=422 n=1024 twiddle= -8.513552e-01   + i -5.245897e-01
		10'd423: twiddle = {-16'd28001   , -16'd17018   }; //i=423 n=1024 twiddle= -8.545580e-01   + i -5.193560e-01
		10'd424: twiddle = {-16'd28105   , -16'd16846   }; //i=424 n=1024 twiddle= -8.577286e-01   + i -5.141027e-01
		10'd425: twiddle = {-16'd28208   , -16'd16673   }; //i=425 n=1024 twiddle= -8.608669e-01   + i -5.088301e-01
		10'd426: twiddle = {-16'd28310   , -16'd16499   }; //i=426 n=1024 twiddle= -8.639729e-01   + i -5.035384e-01
		10'd427: twiddle = {-16'd28411   , -16'd16325   }; //i=427 n=1024 twiddle= -8.670462e-01   + i -4.982277e-01
		10'd428: twiddle = {-16'd28510   , -16'd16151   }; //i=428 n=1024 twiddle= -8.700870e-01   + i -4.928982e-01
		10'd429: twiddle = {-16'd28609   , -16'd15976   }; //i=429 n=1024 twiddle= -8.730950e-01   + i -4.875502e-01
		10'd430: twiddle = {-16'd28706   , -16'd15800   }; //i=430 n=1024 twiddle= -8.760701e-01   + i -4.821838e-01
		10'd431: twiddle = {-16'd28803   , -16'd15623   }; //i=431 n=1024 twiddle= -8.790122e-01   + i -4.767992e-01
		10'd432: twiddle = {-16'd28898   , -16'd15446   }; //i=432 n=1024 twiddle= -8.819213e-01   + i -4.713967e-01
		10'd433: twiddle = {-16'd28992   , -16'd15269   }; //i=433 n=1024 twiddle= -8.847971e-01   + i -4.659765e-01
		10'd434: twiddle = {-16'd29085   , -16'd15090   }; //i=434 n=1024 twiddle= -8.876396e-01   + i -4.605387e-01
		10'd435: twiddle = {-16'd29177   , -16'd14912   }; //i=435 n=1024 twiddle= -8.904487e-01   + i -4.550836e-01
		10'd436: twiddle = {-16'd29268   , -16'd14732   }; //i=436 n=1024 twiddle= -8.932243e-01   + i -4.496113e-01
		10'd437: twiddle = {-16'd29358   , -16'd14553   }; //i=437 n=1024 twiddle= -8.959662e-01   + i -4.441221e-01
		10'd438: twiddle = {-16'd29447   , -16'd14372   }; //i=438 n=1024 twiddle= -8.986745e-01   + i -4.386162e-01
		10'd439: twiddle = {-16'd29534   , -16'd14191   }; //i=439 n=1024 twiddle= -9.013488e-01   + i -4.330938e-01
		10'd440: twiddle = {-16'd29621   , -16'd14010   }; //i=440 n=1024 twiddle= -9.039893e-01   + i -4.275551e-01
		10'd441: twiddle = {-16'd29706   , -16'd13828   }; //i=441 n=1024 twiddle= -9.065957e-01   + i -4.220003e-01
		10'd442: twiddle = {-16'd29791   , -16'd13645   }; //i=442 n=1024 twiddle= -9.091680e-01   + i -4.164296e-01
		10'd443: twiddle = {-16'd29874   , -16'd13462   }; //i=443 n=1024 twiddle= -9.117060e-01   + i -4.108432e-01
		10'd444: twiddle = {-16'd29956   , -16'd13279   }; //i=444 n=1024 twiddle= -9.142098e-01   + i -4.052413e-01
		10'd445: twiddle = {-16'd30037   , -16'd13094   }; //i=445 n=1024 twiddle= -9.166791e-01   + i -3.996242e-01
		10'd446: twiddle = {-16'd30117   , -16'd12910   }; //i=446 n=1024 twiddle= -9.191139e-01   + i -3.939920e-01
		10'd447: twiddle = {-16'd30195   , -16'd12725   }; //i=447 n=1024 twiddle= -9.215140e-01   + i -3.883450e-01
		10'd448: twiddle = {-16'd30273   , -16'd12539   }; //i=448 n=1024 twiddle= -9.238795e-01   + i -3.826834e-01
		10'd449: twiddle = {-16'd30349   , -16'd12353   }; //i=449 n=1024 twiddle= -9.262102e-01   + i -3.770074e-01
		10'd450: twiddle = {-16'd30424   , -16'd12167   }; //i=450 n=1024 twiddle= -9.285061e-01   + i -3.713172e-01
		10'd451: twiddle = {-16'd30498   , -16'd11980   }; //i=451 n=1024 twiddle= -9.307670e-01   + i -3.656130e-01
		10'd452: twiddle = {-16'd30571   , -16'd11793   }; //i=452 n=1024 twiddle= -9.329928e-01   + i -3.598950e-01
		10'd453: twiddle = {-16'd30643   , -16'd11605   }; //i=453 n=1024 twiddle= -9.351835e-01   + i -3.541635e-01
		10'd454: twiddle = {-16'd30714   , -16'd11417   }; //i=454 n=1024 twiddle= -9.373390e-01   + i -3.484187e-01
		10'd455: twiddle = {-16'd30783   , -16'd11228   }; //i=455 n=1024 twiddle= -9.394592e-01   + i -3.426607e-01
		10'd456: twiddle = {-16'd30852   , -16'd11039   }; //i=456 n=1024 twiddle= -9.415441e-01   + i -3.368899e-01
		10'd457: twiddle = {-16'd30919   , -16'd10849   }; //i=457 n=1024 twiddle= -9.435935e-01   + i -3.311063e-01
		10'd458: twiddle = {-16'd30985   , -16'd10659   }; //i=458 n=1024 twiddle= -9.456073e-01   + i -3.253103e-01
		10'd459: twiddle = {-16'd31050   , -16'd10469   }; //i=459 n=1024 twiddle= -9.475856e-01   + i -3.195020e-01
		10'd460: twiddle = {-16'd31113   , -16'd10278   }; //i=460 n=1024 twiddle= -9.495282e-01   + i -3.136817e-01
		10'd461: twiddle = {-16'd31176   , -16'd10087   }; //i=461 n=1024 twiddle= -9.514350e-01   + i -3.078496e-01
		10'd462: twiddle = {-16'd31237   , -16'd9896    }; //i=462 n=1024 twiddle= -9.533060e-01   + i -3.020059e-01
		10'd463: twiddle = {-16'd31297   , -16'd9704    }; //i=463 n=1024 twiddle= -9.551412e-01   + i -2.961509e-01
		10'd464: twiddle = {-16'd31356   , -16'd9512    }; //i=464 n=1024 twiddle= -9.569403e-01   + i -2.902847e-01
		10'd465: twiddle = {-16'd31414   , -16'd9319    }; //i=465 n=1024 twiddle= -9.587035e-01   + i -2.844075e-01
		10'd466: twiddle = {-16'd31470   , -16'd9126    }; //i=466 n=1024 twiddle= -9.604305e-01   + i -2.785197e-01
		10'd467: twiddle = {-16'd31526   , -16'd8933    }; //i=467 n=1024 twiddle= -9.621214e-01   + i -2.726214e-01
		10'd468: twiddle = {-16'd31580   , -16'd8739    }; //i=468 n=1024 twiddle= -9.637761e-01   + i -2.667128e-01
		10'd469: twiddle = {-16'd31633   , -16'd8545    }; //i=469 n=1024 twiddle= -9.653944e-01   + i -2.607941e-01
		10'd470: twiddle = {-16'd31685   , -16'd8351    }; //i=470 n=1024 twiddle= -9.669765e-01   + i -2.548657e-01
		10'd471: twiddle = {-16'd31736   , -16'd8157    }; //i=471 n=1024 twiddle= -9.685221e-01   + i -2.489276e-01
		10'd472: twiddle = {-16'd31785   , -16'd7962    }; //i=472 n=1024 twiddle= -9.700313e-01   + i -2.429802e-01
		10'd473: twiddle = {-16'd31833   , -16'd7767    }; //i=473 n=1024 twiddle= -9.715039e-01   + i -2.370236e-01
		10'd474: twiddle = {-16'd31880   , -16'd7571    }; //i=474 n=1024 twiddle= -9.729400e-01   + i -2.310581e-01
		10'd475: twiddle = {-16'd31926   , -16'd7375    }; //i=475 n=1024 twiddle= -9.743394e-01   + i -2.250839e-01
		10'd476: twiddle = {-16'd31971   , -16'd7179    }; //i=476 n=1024 twiddle= -9.757021e-01   + i -2.191012e-01
		10'd477: twiddle = {-16'd32014   , -16'd6983    }; //i=477 n=1024 twiddle= -9.770281e-01   + i -2.131103e-01
		10'd478: twiddle = {-16'd32057   , -16'd6786    }; //i=478 n=1024 twiddle= -9.783174e-01   + i -2.071114e-01
		10'd479: twiddle = {-16'd32098   , -16'd6590    }; //i=479 n=1024 twiddle= -9.795698e-01   + i -2.011046e-01
		10'd480: twiddle = {-16'd32137   , -16'd6393    }; //i=480 n=1024 twiddle= -9.807853e-01   + i -1.950903e-01
		10'd481: twiddle = {-16'd32176   , -16'd6195    }; //i=481 n=1024 twiddle= -9.819639e-01   + i -1.890687e-01
		10'd482: twiddle = {-16'd32213   , -16'd5998    }; //i=482 n=1024 twiddle= -9.831055e-01   + i -1.830399e-01
		10'd483: twiddle = {-16'd32250   , -16'd5800    }; //i=483 n=1024 twiddle= -9.842101e-01   + i -1.770042e-01
		10'd484: twiddle = {-16'd32285   , -16'd5602    }; //i=484 n=1024 twiddle= -9.852776e-01   + i -1.709619e-01
		10'd485: twiddle = {-16'd32318   , -16'd5404    }; //i=485 n=1024 twiddle= -9.863081e-01   + i -1.649131e-01
		10'd486: twiddle = {-16'd32351   , -16'd5205    }; //i=486 n=1024 twiddle= -9.873014e-01   + i -1.588581e-01
		10'd487: twiddle = {-16'd32382   , -16'd5007    }; //i=487 n=1024 twiddle= -9.882576e-01   + i -1.527972e-01
		10'd488: twiddle = {-16'd32412   , -16'd4808    }; //i=488 n=1024 twiddle= -9.891765e-01   + i -1.467305e-01
		10'd489: twiddle = {-16'd32441   , -16'd4609    }; //i=489 n=1024 twiddle= -9.900582e-01   + i -1.406582e-01
		10'd490: twiddle = {-16'd32469   , -16'd4410    }; //i=490 n=1024 twiddle= -9.909026e-01   + i -1.345807e-01
		10'd491: twiddle = {-16'd32495   , -16'd4210    }; //i=491 n=1024 twiddle= -9.917098e-01   + i -1.284981e-01
		10'd492: twiddle = {-16'd32521   , -16'd4011    }; //i=492 n=1024 twiddle= -9.924795e-01   + i -1.224107e-01
		10'd493: twiddle = {-16'd32545   , -16'd3811    }; //i=493 n=1024 twiddle= -9.932119e-01   + i -1.163186e-01
		10'd494: twiddle = {-16'd32567   , -16'd3612    }; //i=494 n=1024 twiddle= -9.939070e-01   + i -1.102222e-01
		10'd495: twiddle = {-16'd32589   , -16'd3412    }; //i=495 n=1024 twiddle= -9.945646e-01   + i -1.041216e-01
		10'd496: twiddle = {-16'd32609   , -16'd3212    }; //i=496 n=1024 twiddle= -9.951847e-01   + i -9.801714e-02
		10'd497: twiddle = {-16'd32628   , -16'd3012    }; //i=497 n=1024 twiddle= -9.957674e-01   + i -9.190896e-02
		10'd498: twiddle = {-16'd32646   , -16'd2811    }; //i=498 n=1024 twiddle= -9.963126e-01   + i -8.579731e-02
		10'd499: twiddle = {-16'd32663   , -16'd2611    }; //i=499 n=1024 twiddle= -9.968203e-01   + i -7.968244e-02
		10'd500: twiddle = {-16'd32678   , -16'd2410    }; //i=500 n=1024 twiddle= -9.972905e-01   + i -7.356456e-02
		10'd501: twiddle = {-16'd32692   , -16'd2210    }; //i=501 n=1024 twiddle= -9.977231e-01   + i -6.744392e-02
		10'd502: twiddle = {-16'd32705   , -16'd2009    }; //i=502 n=1024 twiddle= -9.981181e-01   + i -6.132074e-02
		10'd503: twiddle = {-16'd32717   , -16'd1809    }; //i=503 n=1024 twiddle= -9.984756e-01   + i -5.519524e-02
		10'd504: twiddle = {-16'd32728   , -16'd1608    }; //i=504 n=1024 twiddle= -9.987955e-01   + i -4.906767e-02
		10'd505: twiddle = {-16'd32737   , -16'd1407    }; //i=505 n=1024 twiddle= -9.990777e-01   + i -4.293826e-02
		10'd506: twiddle = {-16'd32745   , -16'd1206    }; //i=506 n=1024 twiddle= -9.993224e-01   + i -3.680722e-02
		10'd507: twiddle = {-16'd32752   , -16'd1005    }; //i=507 n=1024 twiddle= -9.995294e-01   + i -3.067480e-02
		10'd508: twiddle = {-16'd32757   , -16'd804     }; //i=508 n=1024 twiddle= -9.996988e-01   + i -2.454123e-02
		10'd509: twiddle = {-16'd32761   , -16'd603     }; //i=509 n=1024 twiddle= -9.998306e-01   + i -1.840673e-02
		10'd510: twiddle = {-16'd32765   , -16'd402     }; //i=510 n=1024 twiddle= -9.999247e-01   + i -1.227154e-02
		10'd511: twiddle = {-16'd32766   , -16'd201     }; //i=511 n=1024 twiddle= -9.999812e-01   + i -6.135885e-03
		default: twiddle = 'bX;
		endcase
	end

endmodule