module dualport_ram (
	input Clk, 
	input WE_top, WE_bot,
	input Reset,
	input wire [7:0] addr_top, addr_bot,
	input wire signed [31:0] din_top_re, din_top_im, din_bot_re, din_bot_im,
	output wire signed [31:0] dout_top_re, dout_top_im, dout_bot_re, dout_bot_im
);	

	// RAMB16_S36_S36: 512 x 32 + 4 Parity bits Dual-Port RAM
  //                 Spartan-3E
  // Xilinx HDL Language Template, version 13.1

  RAMB16_S36_S36 #(
     .INIT_A(36'h000000000),  // Value of output RAM registers on Port A at startup
     .INIT_B(36'h000000000),  // Value of output RAM registers on Port B at startup
     .SRVAL_A(36'h000000000), // Port A output value upon SSR assertion
     .SRVAL_B(36'h000000000), // Port B output value upon SSR assertion
     .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
     .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
     .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

     // The following INIT_xx declarations specify the initial contents of the RAM
     // Address 0 to 127
     .INIT_00(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_01(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_02(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_03(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_04(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     // Address 128 to 255
     .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

     // The next set of INITP_xx are for the parity bits
     // Address 0 to 127
     .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
     // Address 128 to 255
     .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) X_Re (
     .DOA(dout_top_re),      // Port A 32-bit Data Output
     .DOB(dout_bot_re),      // Port B 32-bit Data Output
     .DOPA(),    // Port A 4-bit Parity Output
     .DOPB(),    // Port B 4-bit Parity Output
     .ADDRA({1'b1, addr_top}),  // Port A 9-bit Address Input
     .ADDRB({1'b1, addr_bot}),  // Port B 9-bit Address Input
     .CLKA(Clk),    // Port A Clock
     .CLKB(Clk),    // Port B Clock
     .DIA(din_top_re),      // Port A 32-bit Data Input
     .DIB(din_bot_re),      // Port B 32-bit Data Input
     .DIPA(4'd0),    // Port A 4-bit parity Input
     .DIPB(4'd0),    // Port-B 4-bit parity Input
     .ENA(1'b1),      // Port A RAM Enable Input
     .ENB(1'b1),      // Port B RAM Enable Input
     .SSRA(Reset),    // Port A Synchronous Set/Reset Input
     .SSRB(Reset),    // Port B Synchronous Set/Reset Input
     .WEA(WE_top),      // Port A Write Enable Input
     .WEB(WE_bot)       // Port B Write Enable Input
  );
  
  RAMB16_S36_S36 #(
     .INIT_A(36'h000000000),  // Value of output RAM registers on Port A at startup
     .INIT_B(36'h000000000),  // Value of output RAM registers on Port B at startup
     .SRVAL_A(36'h000000000), // Port A output value upon SSR assertion
     .SRVAL_B(36'h000000000), // Port B output value upon SSR assertion
     .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
     .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
     .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

     // The following INIT_xx declarations specify the initial contents of the RAM
     // Address 0 to 127
     .INIT_00(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_01(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_02(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_03(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_04(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     // Address 128 to 255
     .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
     .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

     // The next set of INITP_xx are for the parity bits
     // Address 0 to 127
     .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
     // Address 128 to 255
     .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) X_Im (
     .DOA(dout_top_im),      // Port A 32-bit Data Output
     .DOB(dout_bot_im),      // Port B 32-bit Data Output
     .DOPA(),    // Port A 4-bit Parity Output
     .DOPB(),    // Port B 4-bit Parity Output
     .ADDRA({1'b1, addr_top}),  // Port A 9-bit Address Input
     .ADDRB({1'b1, addr_bot}),  // Port B 9-bit Address Input
     .CLKA(Clk),    // Port A Clock
     .CLKB(Clk),    // Port B Clock
     .DIA(din_top_im),      // Port A 32-bit Data Input
     .DIB(din_bot_im),      // Port B 32-bit Data Input
     .DIPA(4'd0),    // Port A 4-bit parity Input
     .DIPB(4'd0),    // Port-B 4-bit parity Input
     .ENA(1'b1),      // Port A RAM Enable Input
     .ENB(1'b1),      // Port B RAM Enable Input
     .SSRA(Reset),    // Port A Synchronous Set/Reset Input
     .SSRB(Reset),    // Port B Synchronous Set/Reset Input
     .WEA(WE_top),      // Port A Write Enable Input
     .WEB(WE_bot)       // Port B Write Enable Input
  );
  
	

	always@(posedge Clk)
	begin
		$display("-----WE top %b bot %b addr_top %d addr_bot %d data_top_in %d data_top_out %d data_bot_in %d data_bot_out %d", WE_top, WE_bot, addr_top, addr_bot, din_top_re, dout_top_re, din_bot_re, dout_bot_re);
		
	end
    
endmodule