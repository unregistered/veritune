`timescale 1ns / 1ps

module FFT1024_tb_v;
	parameter PRE = 32;
		
	reg Clk;
	reg Reset, Start, Ack;
	reg signed [PRE-1:0] X_Re [1023:0];
	reg signed [PRE-1:0] X_Im [1023:0];
	integer timestamp;
	
	// Outputs
	wire [3:0] state;
	wire Done;
	wire signed [31:0] x_top_re;
	wire signed [31:0] x_top_im;
	wire signed [31:0] x_bot_re;
	wire signed [31:0] x_bot_im;	
	
	// Internal
	wire signed [31:0] y_top_re;
	wire signed [31:0] y_top_im;
	wire signed [31:0] y_bot_re;
	wire signed [31:0] y_bot_im;
	wire [9:0]  i_top, i_bot;
	
	wire signed [31:0] x0, x1, x2, x3, x4, x5, x6, x7;
	assign x0 = X_Re[0];
	assign x1 = X_Re[1];
	assign x2 = X_Re[2];
	assign x3 = X_Re[3];
	assign x4 = X_Re[4];
	assign x5 = X_Re[5];
	assign x6 = X_Re[6];
	assign x7 = X_Re[7];
	assign x_top_re = X_Re[i_top];
	assign x_top_im = X_Im[i_top];
	assign x_bot_re = X_Re[i_bot];
	assign x_bot_im = X_Im[i_bot];
	
	
	// Instantiate the Unit Under Test (UUT)
	FFT1024 uut (
		//	Ins
		.Clk(Clk),
		.Reset(Reset),
		.Start(Start),
		.Ack(Ack),
		.x_top_re(X_Re[i_top]),
		.x_top_im(X_Im[i_top]),
		.x_bot_re(X_Re[i_bot]),
		.x_bot_im(X_Im[i_bot]),
		//	Outs
		.i_top(i_top),
		.i_bot(i_bot),
		.y_top_re(y_top_re),
		.y_top_im(y_top_im),
		.y_bot_re(y_bot_re),
		.y_bot_im(y_bot_im),
		.Done(Done),
		.state(state)
	);
	
	
	initial
	begin
		Clk = 0; // Initialize clock
		Start = 0;
		Reset = 0;
	end
	
	// Keep clock running
	always
	begin
		#20; 
		Clk = ~ Clk; 
	end
	
	//	Here's how to use the butterfly unit
	always @(posedge Clk)
	begin
		timestamp <= timestamp + 1;
		case(state)
			4'd1: //Done
			begin
				$display("X[0]=%d + i%d", X_Re[0], X_Im[0]);
				$display("X[1]=%d + i%d", X_Re[1], X_Im[1]);
				$display("X[2]=%d + i%d", X_Re[2], X_Im[2]);
				$display("X[3]=%d + i%d", X_Re[3], X_Im[3]);
				$display("X[4]=%d + i%d", X_Re[4], X_Im[4]);
				$display("X[5]=%d + i%d", X_Re[5], X_Im[5]);
				$display("X[6]=%d + i%d", X_Re[6], X_Im[6]);
				$display("X[7]=%d + i%d", X_Re[7], X_Im[7]);
				Ack = 1;
			end
			4'd2: //Proc
			begin
				$display("Time: %d", timestamp);
				$display("  i_top %b i_bot %b", i_top, i_bot);
				$display("  x_top_re %d x_bot_re %d", X_Re[i_top], X_Re[i_bot]);
				$display("  y_top %d + i%d y_bot %d + i%d", y_top_re, y_top_im, y_bot_re, y_bot_im);
				X_Re[i_top] <= y_top_re;
				X_Im[i_top] <= y_top_im;
				X_Re[i_bot] <= y_bot_re;
				X_Im[i_bot] <= y_bot_im;
			end
		endcase
	end
	
	//	Just setup
	initial
	begin
		timestamp = 0;
		Start = 0;
		Reset = 0;
		Ack = 0;
		#10
		Reset = 1;
		#200
		// FFT
		X_Re[0]=32'd0;X_Re[512]=-32'd202;X_Re[256]=-32'd2459;X_Re[768]=-32'd1021;X_Re[128]=32'd202;X_Re[640]=32'd1248;X_Re[384]=32'd618;X_Re[896]=-32'd820;X_Re[64]=-32'd1021;X_Re[576]=-32'd2459;X_Re[320]=-32'd4123;X_Re[832]=-32'd4728;X_Re[192]=-32'd5939;X_Re[704]=-32'd6241;X_Re[448]=-32'd2459;X_Re[960]=-32'd416;X_Re[32]=-32'd1248;X_Re[544]=-32'd2459;X_Re[288]=32'd0;X_Re[800]=32'd2459;X_Re[160]=32'd4123;X_Re[672]=32'd5939;X_Re[416]=32'd4930;X_Re[928]=32'd4123;X_Re[96]=32'd2660;X_Re[608]=32'd1853;X_Re[352]=32'd0;X_Re[864]=-32'd2055;X_Re[224]=-32'd3114;X_Re[736]=-32'd1248;X_Re[480]=-32'd202;X_Re[992]=-32'd618;X_Re[16]=-32'd2459;X_Re[528]=-32'd3114;X_Re[272]=-32'd2459;X_Re[784]=-32'd2459;X_Re[144]=-32'd1021;X_Re[656]=-32'd1853;X_Re[400]=-32'd618;X_Re[912]=32'd820;X_Re[80]=32'd1853;X_Re[592]=32'd1853;X_Re[336]=32'd820;X_Re[848]=-32'd618;X_Re[208]=32'd820;X_Re[720]=32'd3518;X_Re[464]=32'd4123;X_Re[976]=32'd2660;X_Re[48]=32'd1021;X_Re[560]=32'd202;X_Re[304]=-32'd1021;X_Re[816]=32'd202;X_Re[176]=-32'd202;X_Re[688]=32'd820;X_Re[432]=32'd3921;X_Re[944]=32'd4930;X_Re[112]=32'd5334;X_Re[624]=32'd5334;X_Re[368]=32'd1652;X_Re[880]=32'd0;X_Re[240]=32'd202;X_Re[752]=-32'd202;X_Re[496]=-32'd3114;X_Re[1008]=-32'd4123;X_Re[8]=-32'd4123;X_Re[520]=-32'd3720;X_Re[264]=-32'd1652;X_Re[776]=-32'd202;X_Re[136]=-32'd618;X_Re[648]=32'd618;X_Re[392]=32'd2660;X_Re[904]=32'd4728;X_Re[72]=32'd4930;X_Re[584]=32'd3518;X_Re[328]=32'd1652;X_Re[840]=32'd1853;X_Re[200]=32'd3921;X_Re[712]=32'd2459;X_Re[456]=32'd820;X_Re[968]=-32'd416;X_Re[40]=32'd618;X_Re[552]=32'd820;X_Re[296]=32'd1853;X_Re[808]=32'd1853;X_Re[168]=32'd1652;X_Re[680]=32'd820;X_Re[424]=-32'd202;X_Re[936]=-32'd820;X_Re[104]=-32'd1652;X_Re[616]=-32'd4728;X_Re[360]=-32'd3316;X_Re[872]=32'd1450;X_Re[232]=32'd2257;X_Re[744]=32'd1021;X_Re[488]=-32'd202;X_Re[1000]=32'd0;X_Re[24]=32'd0;X_Re[536]=32'd2055;X_Re[280]=32'd3114;X_Re[792]=32'd2660;X_Re[152]=32'd3114;X_Re[664]=32'd2257;X_Re[408]=32'd1248;X_Re[920]=32'd618;X_Re[88]=-32'd3114;X_Re[600]=-32'd3518;X_Re[344]=-32'd618;X_Re[856]=32'd1652;X_Re[216]=32'd1652;X_Re[728]=32'd1450;X_Re[472]=32'd416;X_Re[984]=-32'd1853;X_Re[56]=-32'd2257;X_Re[568]=-32'd2459;X_Re[312]=-32'd2660;X_Re[824]=-32'd2459;X_Re[184]=-32'd3518;X_Re[696]=-32'd2913;X_Re[440]=-32'd2257;X_Re[952]=-32'd3316;X_Re[120]=-32'd4930;X_Re[632]=-32'd2459;X_Re[376]=32'd1853;X_Re[888]=32'd2913;X_Re[248]=32'd4123;X_Re[760]=32'd3921;X_Re[504]=32'd1853;X_Re[1016]=32'd820;X_Re[4]=32'd2257;X_Re[516]=32'd1652;X_Re[260]=32'd820;X_Re[772]=32'd618;X_Re[132]=32'd1021;X_Re[644]=32'd1652;X_Re[388]=32'd416;X_Re[900]=-32'd2055;X_Re[68]=-32'd2660;X_Re[580]=-32'd2660;X_Re[324]=-32'd3518;X_Re[836]=-32'd3114;X_Re[196]=-32'd3518;X_Re[708]=-32'd3518;X_Re[452]=-32'd3114;X_Re[964]=-32'd202;X_Re[36]=32'd202;X_Re[548]=32'd416;X_Re[292]=32'd1853;X_Re[804]=32'd1853;X_Re[164]=32'd1853;X_Re[676]=32'd2257;X_Re[420]=32'd820;X_Re[932]=-32'd820;X_Re[100]=32'd618;X_Re[612]=32'd1248;X_Re[356]=32'd820;X_Re[868]=-32'd202;X_Re[228]=-32'd618;X_Re[740]=-32'd618;X_Re[484]=32'd1021;X_Re[996]=32'd3114;X_Re[20]=32'd3114;X_Re[532]=32'd3720;X_Re[276]=32'd1248;X_Re[788]=-32'd416;X_Re[148]=-32'd1652;X_Re[660]=-32'd5132;X_Re[404]=-32'd7452;X_Re[916]=-32'd6241;X_Re[84]=-32'd3720;X_Re[596]=-32'd2257;X_Re[340]=-32'd202;X_Re[852]=32'd202;X_Re[212]=-32'd416;X_Re[724]=32'd1450;X_Re[468]=32'd3921;X_Re[980]=32'd4325;X_Re[52]=32'd4930;X_Re[564]=32'd5132;X_Re[308]=32'd4123;X_Re[820]=32'd3518;X_Re[180]=32'd1248;X_Re[692]=-32'd1652;X_Re[436]=-32'd3518;X_Re[948]=-32'd1652;X_Re[116]=32'd618;X_Re[628]=32'd1021;X_Re[372]=32'd1652;X_Re[884]=32'd0;X_Re[244]=-32'd1248;X_Re[756]=-32'd1450;X_Re[500]=-32'd2055;X_Re[1012]=-32'd1450;X_Re[12]=-32'd202;X_Re[524]=32'd0;X_Re[268]=32'd416;X_Re[780]=32'd820;X_Re[140]=-32'd618;X_Re[652]=-32'd1652;X_Re[396]=-32'd618;X_Re[908]=32'd1021;X_Re[76]=32'd1652;X_Re[588]=32'd3720;X_Re[332]=32'd2913;X_Re[844]=32'd1248;X_Re[204]=32'd1021;X_Re[716]=32'd1450;X_Re[460]=32'd1021;X_Re[972]=32'd820;X_Re[44]=32'd1450;X_Re[556]=32'd1853;X_Re[300]=32'd2660;X_Re[812]=32'd2055;X_Re[172]=32'd1021;X_Re[684]=-32'd202;X_Re[428]=-32'd416;X_Re[940]=-32'd618;X_Re[108]=-32'd416;X_Re[620]=-32'd1853;X_Re[364]=-32'd3921;X_Re[876]=-32'd4123;X_Re[236]=-32'd3921;X_Re[748]=-32'd3921;X_Re[492]=-32'd2459;X_Re[1004]=-32'd1021;X_Re[28]=-32'd1450;X_Re[540]=-32'd416;X_Re[284]=32'd618;X_Re[796]=32'd618;X_Re[156]=32'd1021;X_Re[668]=32'd2660;X_Re[412]=32'd4527;X_Re[924]=32'd4728;X_Re[92]=32'd4123;X_Re[604]=32'd416;X_Re[348]=-32'd820;X_Re[860]=-32'd416;X_Re[220]=32'd416;X_Re[732]=32'd202;X_Re[476]=32'd1021;X_Re[988]=32'd202;X_Re[60]=-32'd1853;X_Re[572]=-32'd4325;X_Re[316]=-32'd5334;X_Re[828]=-32'd5535;X_Re[188]=-32'd4728;X_Re[700]=-32'd2660;X_Re[444]=-32'd202;X_Re[956]=32'd1450;X_Re[124]=32'd1450;X_Re[636]=32'd1021;X_Re[380]=32'd1652;X_Re[892]=32'd1248;X_Re[252]=32'd1021;X_Re[764]=32'd2257;X_Re[508]=32'd2660;X_Re[1020]=32'd820;X_Re[2]=32'd0;X_Re[514]=-32'd1021;X_Re[258]=-32'd3114;X_Re[770]=-32'd3316;X_Re[130]=32'd416;X_Re[642]=32'd2459;X_Re[386]=32'd4123;X_Re[898]=32'd3921;X_Re[66]=32'd2459;X_Re[578]=32'd1248;X_Re[322]=32'd0;X_Re[834]=-32'd1652;X_Re[194]=-32'd2257;X_Re[706]=-32'd2257;X_Re[450]=-32'd3114;X_Re[962]=-32'd3720;X_Re[34]=-32'd3518;X_Re[546]=-32'd3921;X_Re[290]=-32'd3720;X_Re[802]=-32'd1450;X_Re[162]=32'd1021;X_Re[674]=32'd3720;X_Re[418]=32'd4728;X_Re[930]=32'd3720;X_Re[98]=32'd3316;X_Re[610]=32'd4123;X_Re[354]=32'd3316;X_Re[866]=32'd3114;X_Re[226]=32'd2913;X_Re[738]=32'd1248;X_Re[482]=32'd618;X_Re[994]=32'd820;X_Re[18]=32'd820;X_Re[530]=-32'd618;X_Re[274]=-32'd1021;X_Re[786]=-32'd618;X_Re[146]=-32'd416;X_Re[658]=32'd202;X_Re[402]=-32'd416;X_Re[914]=-32'd1450;X_Re[82]=-32'd2055;X_Re[594]=-32'd1853;X_Re[338]=-32'd1248;X_Re[850]=32'd618;X_Re[210]=32'd820;X_Re[722]=32'd820;X_Re[466]=-32'd416;X_Re[978]=-32'd202;X_Re[50]=-32'd820;X_Re[562]=-32'd202;X_Re[306]=32'd1652;X_Re[818]=32'd3114;X_Re[178]=32'd3921;X_Re[690]=32'd2660;X_Re[434]=32'd202;X_Re[946]=-32'd416;X_Re[114]=32'd1021;X_Re[626]=32'd1021;X_Re[370]=32'd1021;X_Re[882]=32'd3114;X_Re[242]=32'd2257;X_Re[754]=-32'd202;X_Re[498]=-32'd1248;X_Re[1010]=-32'd2660;X_Re[10]=-32'd4728;X_Re[522]=-32'd4325;X_Re[266]=-32'd2660;X_Re[778]=-32'd1450;X_Re[138]=-32'd1652;X_Re[650]=-32'd1248;X_Re[394]=-32'd1021;X_Re[906]=-32'd202;X_Re[74]=-32'd820;X_Re[586]=32'd416;X_Re[330]=32'd1652;X_Re[842]=32'd1853;X_Re[202]=32'd2055;X_Re[714]=32'd1853;X_Re[458]=32'd0;X_Re[970]=-32'd2660;X_Re[42]=-32'd2913;X_Re[554]=-32'd1021;X_Re[298]=32'd1248;X_Re[810]=32'd1450;X_Re[170]=32'd820;X_Re[682]=32'd202;X_Re[426]=-32'd1021;X_Re[938]=-32'd2913;X_Re[106]=-32'd2660;X_Re[618]=-32'd1853;X_Re[362]=-32'd1450;X_Re[874]=-32'd2257;X_Re[234]=-32'd2660;X_Re[746]=-32'd3114;X_Re[490]=-32'd3518;X_Re[1002]=-32'd2660;X_Re[26]=32'd0;X_Re[538]=32'd1652;X_Re[282]=32'd2257;X_Re[794]=32'd1652;X_Re[154]=32'd1021;X_Re[666]=32'd1450;X_Re[410]=32'd1450;X_Re[922]=32'd1021;X_Re[90]=32'd618;X_Re[602]=32'd618;X_Re[346]=32'd416;X_Re[858]=32'd1021;X_Re[218]=32'd2055;X_Re[730]=32'd1021;X_Re[474]=32'd618;X_Re[986]=32'd2257;X_Re[58]=32'd3114;X_Re[570]=32'd3518;X_Re[314]=32'd1853;X_Re[826]=-32'd202;X_Re[186]=-32'd1853;X_Re[698]=-32'd3316;X_Re[442]=-32'd4728;X_Re[954]=-32'd4123;X_Re[122]=-32'd2913;X_Re[634]=-32'd1853;X_Re[378]=-32'd2257;X_Re[890]=-32'd2257;X_Re[250]=-32'd1450;X_Re[762]=-32'd1248;X_Re[506]=32'd820;X_Re[1018]=32'd4527;X_Re[6]=32'd7452;X_Re[518]=32'd7048;X_Re[262]=32'd5132;X_Re[774]=32'd3316;X_Re[134]=32'd1853;X_Re[646]=32'd1021;X_Re[390]=32'd820;X_Re[902]=32'd1450;X_Re[70]=32'd1248;X_Re[582]=-32'd1450;X_Re[326]=-32'd2257;X_Re[838]=-32'd2660;X_Re[198]=-32'd4325;X_Re[710]=-32'd3921;X_Re[454]=-32'd1853;X_Re[966]=32'd618;X_Re[38]=32'd0;X_Re[550]=32'd820;X_Re[294]=32'd2055;X_Re[806]=32'd2055;X_Re[166]=32'd1450;X_Re[678]=32'd1248;X_Re[422]=32'd1450;X_Re[934]=32'd1652;X_Re[102]=32'd618;X_Re[614]=32'd1248;X_Re[358]=32'd820;X_Re[870]=-32'd1652;X_Re[230]=-32'd2257;X_Re[742]=32'd202;X_Re[486]=32'd3114;X_Re[998]=32'd3921;X_Re[22]=32'd3720;X_Re[534]=32'd3518;X_Re[278]=32'd2257;X_Re[790]=32'd820;X_Re[150]=-32'd416;X_Re[662]=-32'd618;X_Re[406]=-32'd820;X_Re[918]=-32'd2055;X_Re[86]=-32'd2660;X_Re[598]=-32'd3316;X_Re[342]=-32'd4930;X_Re[854]=-32'd4930;X_Re[214]=-32'd2459;X_Re[726]=-32'd618;X_Re[470]=32'd1248;X_Re[982]=32'd820;X_Re[54]=32'd2459;X_Re[566]=32'd3114;X_Re[310]=32'd2913;X_Re[822]=32'd2459;X_Re[182]=32'd2459;X_Re[694]=32'd1450;X_Re[438]=32'd1021;X_Re[950]=32'd0;X_Re[118]=-32'd202;X_Re[630]=-32'd618;X_Re[374]=-32'd416;X_Re[886]=32'd416;X_Re[246]=32'd1652;X_Re[758]=32'd2660;X_Re[502]=32'd1450;X_Re[1014]=32'd618;X_Re[14]=32'd0;X_Re[526]=-32'd416;X_Re[270]=-32'd1652;X_Re[782]=-32'd3720;X_Re[142]=-32'd3921;X_Re[654]=-32'd2913;X_Re[398]=-32'd3114;X_Re[910]=-32'd2459;X_Re[78]=-32'd2055;X_Re[590]=-32'd2913;X_Re[334]=-32'd2257;X_Re[846]=32'd1021;X_Re[206]=32'd4325;X_Re[718]=32'd4527;X_Re[462]=32'd2913;X_Re[974]=32'd2055;X_Re[46]=32'd1652;X_Re[558]=32'd618;X_Re[302]=-32'd202;X_Re[814]=32'd1450;X_Re[174]=32'd1853;X_Re[686]=32'd416;X_Re[430]=-32'd820;X_Re[942]=-32'd202;X_Re[110]=-32'd2055;X_Re[622]=-32'd3114;X_Re[366]=-32'd2055;X_Re[878]=-32'd416;X_Re[238]=-32'd618;X_Re[750]=-32'd1652;X_Re[494]=-32'd1248;X_Re[1006]=-32'd1450;X_Re[30]=-32'd2257;X_Re[542]=-32'd2660;X_Re[286]=-32'd1853;X_Re[798]=-32'd1450;X_Re[158]=-32'd1021;X_Re[670]=-32'd416;X_Re[414]=32'd820;X_Re[926]=32'd416;X_Re[94]=-32'd820;X_Re[606]=32'd618;X_Re[350]=32'd2660;X_Re[862]=32'd3316;X_Re[222]=32'd2913;X_Re[734]=32'd2913;X_Re[478]=32'd2055;X_Re[990]=32'd416;X_Re[62]=-32'd1021;X_Re[574]=-32'd1853;X_Re[318]=-32'd1853;X_Re[830]=-32'd1853;X_Re[190]=-32'd2055;X_Re[702]=-32'd1450;X_Re[446]=-32'd1853;X_Re[958]=-32'd3114;X_Re[126]=-32'd1853;X_Re[638]=-32'd202;X_Re[382]=32'd1450;X_Re[894]=32'd1450;X_Re[254]=32'd416;X_Re[766]=32'd416;X_Re[510]=32'd416;X_Re[1022]=32'd618;X_Re[1]=32'd202;X_Re[513]=-32'd202;X_Re[257]=-32'd202;X_Re[769]=32'd0;X_Re[129]=-32'd202;X_Re[641]=32'd416;X_Re[385]=32'd618;X_Re[897]=32'd1853;X_Re[65]=32'd3921;X_Re[577]=32'd5334;X_Re[321]=32'd4527;X_Re[833]=32'd3720;X_Re[193]=32'd2660;X_Re[705]=32'd1450;X_Re[449]=-32'd618;X_Re[961]=-32'd2257;X_Re[33]=-32'd4123;X_Re[545]=-32'd4123;X_Re[289]=-32'd4527;X_Re[801]=-32'd4527;X_Re[161]=-32'd3720;X_Re[673]=-32'd2459;X_Re[417]=-32'd1652;X_Re[929]=32'd1652;X_Re[97]=32'd3921;X_Re[609]=32'd6241;X_Re[353]=32'd5535;X_Re[865]=32'd4728;X_Re[225]=32'd4527;X_Re[737]=32'd3921;X_Re[481]=32'd2257;X_Re[993]=32'd1021;X_Re[17]=32'd820;X_Re[529]=32'd0;X_Re[273]=-32'd820;X_Re[785]=-32'd820;X_Re[145]=-32'd1450;X_Re[657]=-32'd2055;X_Re[401]=-32'd1248;X_Re[913]=32'd1248;X_Re[81]=32'd2660;X_Re[593]=32'd1450;X_Re[337]=32'd1248;X_Re[849]=32'd820;X_Re[209]=32'd618;X_Re[721]=32'd0;X_Re[465]=-32'd202;X_Re[977]=-32'd618;X_Re[49]=-32'd1021;X_Re[561]=-32'd1248;X_Re[305]=-32'd618;X_Re[817]=-32'd202;X_Re[177]=-32'd416;X_Re[689]=-32'd618;X_Re[433]=32'd1021;X_Re[945]=32'd1853;X_Re[113]=32'd2055;X_Re[625]=32'd2257;X_Re[369]=32'd2257;X_Re[881]=32'd2055;X_Re[241]=32'd1248;X_Re[753]=-32'd202;X_Re[497]=-32'd1450;X_Re[1009]=-32'd1652;X_Re[9]=-32'd2055;X_Re[521]=-32'd2660;X_Re[265]=-32'd2913;X_Re[777]=-32'd3114;X_Re[137]=-32'd3316;X_Re[649]=-32'd2660;X_Re[393]=-32'd618;X_Re[905]=-32'd416;X_Re[73]=-32'd618;X_Re[585]=32'd0;X_Re[329]=32'd820;X_Re[841]=32'd1450;X_Re[201]=32'd1450;X_Re[713]=32'd1248;X_Re[457]=32'd0;X_Re[969]=32'd0;X_Re[41]=-32'd618;X_Re[553]=-32'd820;X_Re[297]=-32'd820;X_Re[809]=-32'd1021;X_Re[169]=32'd202;X_Re[681]=32'd1652;X_Re[425]=32'd2257;X_Re[937]=32'd1450;X_Re[105]=32'd618;X_Re[617]=32'd1021;X_Re[361]=32'd1021;X_Re[873]=32'd202;X_Re[233]=-32'd1021;X_Re[745]=-32'd2257;X_Re[489]=-32'd2913;X_Re[1001]=-32'd3316;X_Re[25]=-32'd2459;X_Re[537]=-32'd2660;X_Re[281]=-32'd2459;X_Re[793]=-32'd1652;X_Re[153]=-32'd416;X_Re[665]=32'd1450;X_Re[409]=32'd2055;X_Re[921]=32'd1853;X_Re[89]=32'd2257;X_Re[601]=32'd2660;X_Re[345]=32'd1853;X_Re[857]=32'd820;X_Re[217]=32'd202;X_Re[729]=32'd0;X_Re[473]=-32'd202;X_Re[985]=-32'd202;X_Re[57]=32'd0;X_Re[569]=-32'd618;X_Re[313]=-32'd618;X_Re[825]=32'd820;X_Re[185]=32'd1652;X_Re[697]=32'd1450;X_Re[441]=32'd618;X_Re[953]=-32'd618;X_Re[121]=-32'd1021;X_Re[633]=-32'd1248;X_Re[377]=-32'd1450;X_Re[889]=-32'd2913;X_Re[249]=-32'd3720;X_Re[761]=-32'd2913;X_Re[505]=-32'd1853;X_Re[1017]=-32'd618;X_Re[5]=32'd820;X_Re[517]=32'd1021;X_Re[261]=32'd2257;X_Re[773]=32'd3114;X_Re[133]=32'd3114;X_Re[645]=32'd2459;X_Re[389]=32'd2055;X_Re[901]=32'd1853;X_Re[69]=32'd1450;X_Re[581]=32'd1021;X_Re[325]=32'd0;X_Re[837]=-32'd1652;X_Re[197]=-32'd2055;X_Re[709]=-32'd1450;X_Re[453]=-32'd1021;X_Re[965]=-32'd1021;X_Re[37]=-32'd618;X_Re[549]=-32'd416;X_Re[293]=-32'd416;X_Re[805]=32'd618;X_Re[165]=32'd1248;X_Re[677]=32'd820;X_Re[421]=32'd1450;X_Re[933]=32'd1021;X_Re[101]=32'd618;X_Re[613]=32'd202;X_Re[357]=-32'd202;X_Re[869]=-32'd1021;X_Re[229]=-32'd416;X_Re[741]=-32'd202;X_Re[485]=-32'd416;X_Re[997]=32'd618;X_Re[21]=32'd2257;X_Re[533]=32'd3720;X_Re[277]=32'd4527;X_Re[789]=32'd5132;X_Re[149]=32'd4325;X_Re[661]=32'd3921;X_Re[405]=32'd3720;X_Re[917]=32'd2660;X_Re[85]=32'd202;X_Re[597]=-32'd2055;X_Re[341]=-32'd4325;X_Re[853]=-32'd5132;X_Re[213]=-32'd5535;X_Re[725]=-32'd4930;X_Re[469]=-32'd4325;X_Re[981]=-32'd3720;X_Re[53]=-32'd2055;X_Re[565]=-32'd416;X_Re[309]=32'd1021;X_Re[821]=32'd1853;X_Re[181]=32'd2459;X_Re[693]=32'd3720;X_Re[437]=32'd4728;X_Re[949]=32'd3518;X_Re[117]=32'd2257;X_Re[629]=-32'd202;X_Re[373]=-32'd1248;X_Re[885]=-32'd2257;X_Re[245]=-32'd2257;X_Re[757]=-32'd2660;X_Re[501]=-32'd2257;X_Re[1013]=-32'd1652;X_Re[13]=-32'd202;X_Re[525]=32'd618;X_Re[269]=32'd820;X_Re[781]=32'd618;X_Re[141]=32'd1248;X_Re[653]=32'd1248;X_Re[397]=32'd202;X_Re[909]=-32'd618;X_Re[77]=-32'd2459;X_Re[589]=-32'd3316;X_Re[333]=-32'd3316;X_Re[845]=-32'd3114;X_Re[205]=-32'd2913;X_Re[717]=-32'd1652;X_Re[461]=-32'd618;X_Re[973]=32'd820;X_Re[45]=32'd2055;X_Re[557]=32'd2459;X_Re[301]=32'd2055;X_Re[813]=32'd2055;X_Re[173]=32'd2660;X_Re[685]=32'd2913;X_Re[429]=32'd2257;X_Re[941]=32'd1021;X_Re[109]=-32'd618;X_Re[621]=-32'd820;X_Re[365]=-32'd820;X_Re[877]=-32'd1021;X_Re[237]=-32'd820;X_Re[749]=-32'd416;X_Re[493]=-32'd1021;X_Re[1005]=-32'd1248;X_Re[29]=-32'd1248;X_Re[541]=-32'd618;X_Re[285]=-32'd416;X_Re[797]=32'd202;X_Re[157]=32'd1021;X_Re[669]=32'd1021;X_Re[413]=-32'd202;X_Re[925]=-32'd820;X_Re[93]=32'd0;X_Re[605]=32'd202;X_Re[349]=32'd820;X_Re[861]=32'd820;X_Re[221]=32'd1450;X_Re[733]=32'd1021;X_Re[477]=32'd1450;X_Re[989]=32'd2055;X_Re[61]=32'd2257;X_Re[573]=32'd2913;X_Re[317]=32'd3316;X_Re[829]=32'd3518;X_Re[189]=32'd2459;X_Re[701]=32'd618;X_Re[445]=-32'd820;X_Re[957]=-32'd2459;X_Re[125]=-32'd3114;X_Re[637]=-32'd3316;X_Re[381]=-32'd2913;X_Re[893]=-32'd1853;X_Re[253]=-32'd416;X_Re[765]=32'd202;X_Re[509]=32'd416;X_Re[1021]=32'd618;X_Re[3]=32'd618;X_Re[515]=32'd1853;X_Re[259]=32'd3316;X_Re[771]=32'd3518;X_Re[131]=32'd2913;X_Re[643]=32'd618;X_Re[387]=-32'd1248;X_Re[899]=-32'd1450;X_Re[67]=-32'd820;X_Re[579]=-32'd820;X_Re[323]=-32'd416;X_Re[835]=32'd1021;X_Re[195]=32'd1450;X_Re[707]=32'd1853;X_Re[451]=32'd2055;X_Re[963]=32'd1652;X_Re[35]=32'd1450;X_Re[547]=32'd1248;X_Re[291]=32'd202;X_Re[803]=-32'd1021;X_Re[163]=-32'd2459;X_Re[675]=-32'd3316;X_Re[419]=-32'd3518;X_Re[931]=-32'd2913;X_Re[99]=-32'd2459;X_Re[611]=-32'd2055;X_Re[355]=-32'd1450;X_Re[867]=32'd0;X_Re[227]=32'd1021;X_Re[739]=32'd2055;X_Re[483]=32'd2660;X_Re[995]=32'd2257;X_Re[19]=32'd1450;X_Re[531]=32'd1652;X_Re[275]=32'd1021;X_Re[787]=-32'd820;X_Re[147]=-32'd2660;X_Re[659]=-32'd2660;X_Re[403]=-32'd3114;X_Re[915]=-32'd2257;X_Re[83]=-32'd1652;X_Re[595]=-32'd1021;X_Re[339]=32'd202;X_Re[851]=32'd416;X_Re[211]=-32'd202;X_Re[723]=32'd202;X_Re[467]=32'd416;X_Re[979]=32'd416;X_Re[51]=32'd820;X_Re[563]=32'd618;X_Re[307]=-32'd1021;X_Re[819]=-32'd3114;X_Re[179]=-32'd3518;X_Re[691]=-32'd3518;X_Re[435]=-32'd1853;X_Re[947]=-32'd618;X_Re[115]=32'd618;X_Re[627]=32'd1021;X_Re[371]=32'd1450;X_Re[883]=32'd1853;X_Re[243]=32'd2055;X_Re[755]=32'd2055;X_Re[499]=32'd2459;X_Re[1011]=32'd3316;X_Re[11]=32'd3316;X_Re[523]=32'd2459;X_Re[267]=32'd1021;X_Re[779]=-32'd1021;X_Re[139]=-32'd2055;X_Re[651]=-32'd2660;X_Re[395]=-32'd3518;X_Re[907]=-32'd3316;X_Re[75]=-32'd1652;X_Re[587]=-32'd202;X_Re[331]=32'd202;X_Re[843]=32'd416;X_Re[203]=32'd1021;X_Re[715]=32'd1652;X_Re[459]=32'd2660;X_Re[971]=32'd3316;X_Re[43]=32'd4527;X_Re[555]=32'd3316;X_Re[299]=32'd1450;X_Re[811]=-32'd202;X_Re[171]=-32'd1652;X_Re[683]=-32'd1450;X_Re[427]=-32'd1853;X_Re[939]=-32'd1248;X_Re[107]=32'd0;X_Re[619]=32'd1021;X_Re[363]=32'd1248;X_Re[875]=32'd2660;X_Re[235]=32'd2660;X_Re[747]=32'd2660;X_Re[491]=32'd3518;X_Re[1003]=32'd2257;X_Re[27]=-32'd202;X_Re[539]=-32'd1652;X_Re[283]=-32'd2055;X_Re[795]=-32'd2257;X_Re[155]=-32'd1652;X_Re[667]=-32'd1652;X_Re[411]=-32'd1450;X_Re[923]=-32'd1021;X_Re[91]=-32'd820;X_Re[603]=-32'd820;X_Re[347]=32'd202;X_Re[859]=32'd1450;X_Re[219]=32'd1248;X_Re[731]=32'd1853;X_Re[475]=32'd2459;X_Re[987]=32'd1853;X_Re[59]=-32'd202;X_Re[571]=-32'd202;X_Re[315]=-32'd820;X_Re[827]=-32'd618;X_Re[187]=32'd416;X_Re[699]=32'd1021;X_Re[443]=32'd416;X_Re[955]=32'd820;X_Re[123]=32'd416;X_Re[635]=-32'd618;X_Re[379]=-32'd416;X_Re[891]=-32'd202;X_Re[251]=32'd416;X_Re[763]=32'd820;X_Re[507]=32'd618;X_Re[1019]=-32'd1652;X_Re[7]=-32'd2459;X_Re[519]=-32'd3114;X_Re[263]=-32'd3114;X_Re[775]=-32'd1248;X_Re[135]=32'd1021;X_Re[647]=32'd1248;X_Re[391]=32'd2257;X_Re[903]=32'd2913;X_Re[71]=32'd2055;X_Re[583]=32'd2257;X_Re[327]=32'd2660;X_Re[839]=32'd2257;X_Re[199]=32'd2660;X_Re[711]=32'd3114;X_Re[455]=32'd1652;X_Re[967]=-32'd416;X_Re[39]=-32'd1450;X_Re[551]=-32'd2055;X_Re[295]=-32'd2913;X_Re[807]=-32'd2660;X_Re[167]=-32'd2913;X_Re[679]=-32'd2055;X_Re[423]=-32'd1450;X_Re[935]=-32'd1248;X_Re[103]=-32'd1021;X_Re[615]=-32'd416;X_Re[359]=-32'd202;X_Re[871]=32'd0;X_Re[231]=32'd820;X_Re[743]=32'd820;X_Re[487]=32'd202;X_Re[999]=32'd0;X_Re[23]=-32'd618;X_Re[535]=-32'd820;X_Re[279]=-32'd1248;X_Re[791]=-32'd1248;X_Re[151]=-32'd1021;X_Re[663]=-32'd202;X_Re[407]=32'd618;X_Re[919]=32'd1450;X_Re[87]=32'd2257;X_Re[599]=32'd2660;X_Re[343]=32'd2913;X_Re[855]=32'd2660;X_Re[215]=32'd1021;X_Re[727]=-32'd1021;X_Re[471]=-32'd3114;X_Re[983]=-32'd3720;X_Re[55]=-32'd3518;X_Re[567]=-32'd3518;X_Re[311]=-32'd2055;X_Re[823]=-32'd1853;X_Re[183]=-32'd202;X_Re[695]=32'd0;X_Re[439]=32'd0;X_Re[951]=32'd1248;X_Re[119]=32'd2257;X_Re[631]=32'd2660;X_Re[375]=32'd3720;X_Re[887]=32'd3720;X_Re[247]=32'd1450;X_Re[759]=-32'd618;X_Re[503]=-32'd1652;X_Re[1015]=-32'd2459;X_Re[15]=-32'd1853;X_Re[527]=-32'd618;X_Re[271]=-32'd820;X_Re[783]=32'd618;X_Re[143]=32'd1652;X_Re[655]=32'd1021;X_Re[399]=32'd416;X_Re[911]=32'd618;X_Re[79]=32'd618;X_Re[591]=32'd820;X_Re[335]=32'd1652;X_Re[847]=32'd416;X_Re[207]=-32'd1021;X_Re[719]=-32'd2913;X_Re[463]=-32'd3114;X_Re[975]=-32'd3518;X_Re[47]=-32'd2913;X_Re[559]=-32'd1853;X_Re[303]=-32'd416;X_Re[815]=32'd1021;X_Re[175]=32'd1652;X_Re[687]=32'd1853;X_Re[431]=32'd2660;X_Re[943]=32'd2459;X_Re[111]=32'd2055;X_Re[623]=32'd2913;X_Re[367]=32'd2913;X_Re[879]=32'd618;X_Re[239]=-32'd1021;X_Re[751]=-32'd1248;X_Re[495]=-32'd1853;X_Re[1007]=-32'd1853;X_Re[31]=-32'd1652;X_Re[543]=-32'd2257;X_Re[287]=-32'd1450;X_Re[799]=-32'd416;X_Re[159]=32'd0;X_Re[671]=32'd1248;X_Re[415]=32'd1853;X_Re[927]=32'd2055;X_Re[95]=32'd2660;X_Re[607]=32'd2055;X_Re[351]=32'd820;X_Re[863]=-32'd416;X_Re[223]=-32'd1450;X_Re[735]=-32'd1021;X_Re[479]=-32'd1021;X_Re[991]=-32'd618;X_Re[63]=-32'd820;X_Re[575]=-32'd618;X_Re[319]=-32'd202;X_Re[831]=32'd202;X_Re[191]=32'd1021;X_Re[703]=32'd1853;X_Re[447]=32'd3114;X_Re[959]=32'd3921;X_Re[127]=32'd4123;X_Re[639]=32'd2660;X_Re[383]=32'd416;X_Re[895]=-32'd1248;X_Re[255]=-32'd1450;X_Re[767]=-32'd1652;X_Re[511]=-32'd1450;X_Re[1023]=-32'd1450;
		X_Im[0]=32'd0; X_Im[1]=-32'd0; X_Im[2]=-32'd0; X_Im[3]=-32'd0; X_Im[4]=32'd0; X_Im[5]=32'd0; X_Im[6]=32'd0; X_Im[7]=-32'd0; X_Im[8]=-32'd0; X_Im[9]=-32'd0; X_Im[10]=-32'd0; X_Im[11]=-32'd0; X_Im[12]=-32'd0; X_Im[13]=-32'd0; X_Im[14]=-32'd0; X_Im[15]=-32'd0; X_Im[16]=-32'd0; X_Im[17]=-32'd0; X_Im[18]=32'd0; X_Im[19]=32'd0; X_Im[20]=32'd0; X_Im[21]=32'd0; X_Im[22]=32'd0; X_Im[23]=32'd0; X_Im[24]=32'd0; X_Im[25]=32'd0; X_Im[26]=32'd0; X_Im[27]=-32'd0; X_Im[28]=-32'd0; X_Im[29]=-32'd0; X_Im[30]=-32'd0; X_Im[31]=-32'd0; X_Im[32]=-32'd0; X_Im[33]=-32'd0; X_Im[34]=-32'd0; X_Im[35]=-32'd0; X_Im[36]=-32'd0; X_Im[37]=-32'd0; X_Im[38]=-32'd0; X_Im[39]=32'd0; X_Im[40]=32'd0; X_Im[41]=32'd0; X_Im[42]=32'd0; X_Im[43]=-32'd0; X_Im[44]=32'd0; X_Im[45]=32'd0; X_Im[46]=32'd0; X_Im[47]=32'd0; X_Im[48]=32'd0; X_Im[49]=32'd0; X_Im[50]=-32'd0; X_Im[51]=32'd0; X_Im[52]=-32'd0; X_Im[53]=32'd0; X_Im[54]=32'd0; X_Im[55]=32'd0; X_Im[56]=32'd0; X_Im[57]=32'd0; X_Im[58]=32'd0; X_Im[59]=32'd0; X_Im[60]=32'd0; X_Im[61]=-32'd0; X_Im[62]=-32'd0; X_Im[63]=-32'd0; X_Im[64]=-32'd0; X_Im[65]=-32'd0; X_Im[66]=-32'd0; X_Im[67]=-32'd0; X_Im[68]=-32'd0; X_Im[69]=32'd0; X_Im[70]=32'd0; X_Im[71]=32'd0; X_Im[72]=32'd0; X_Im[73]=32'd0; X_Im[74]=32'd0; X_Im[75]=32'd0; X_Im[76]=32'd0; X_Im[77]=32'd0; X_Im[78]=32'd0; X_Im[79]=-32'd0; X_Im[80]=32'd0; X_Im[81]=32'd0; X_Im[82]=32'd0; X_Im[83]=32'd0; X_Im[84]=32'd0; X_Im[85]=32'd0; X_Im[86]=-32'd0; X_Im[87]=-32'd0; X_Im[88]=-32'd0; X_Im[89]=-32'd0; X_Im[90]=-32'd0; X_Im[91]=32'd0; X_Im[92]=32'd0; X_Im[93]=32'd0; X_Im[94]=-32'd0; X_Im[95]=32'd0; X_Im[96]=32'd0; X_Im[97]=32'd0; X_Im[98]=32'd0; X_Im[99]=32'd0; X_Im[100]=32'd0; X_Im[101]=32'd0; X_Im[102]=32'd0; X_Im[103]=32'd0; X_Im[104]=-32'd0; X_Im[105]=-32'd0; X_Im[106]=-32'd0; X_Im[107]=32'd0; X_Im[108]=32'd0; X_Im[109]=32'd0; X_Im[110]=32'd0; X_Im[111]=-32'd0; X_Im[112]=-32'd0; X_Im[113]=-32'd0; X_Im[114]=-32'd0; X_Im[115]=-32'd0; X_Im[116]=-32'd0; X_Im[117]=-32'd0; X_Im[118]=-32'd0; X_Im[119]=-32'd0; X_Im[120]=-32'd0; X_Im[121]=-32'd0; X_Im[122]=32'd0; X_Im[123]=32'd0; X_Im[124]=32'd0; X_Im[125]=32'd0; X_Im[126]=32'd0; X_Im[127]=32'd0; X_Im[128]=32'd0; X_Im[129]=32'd0; X_Im[130]=32'd0; X_Im[131]=32'd0; X_Im[132]=32'd0; X_Im[133]=32'd0; X_Im[134]=32'd0; X_Im[135]=-32'd0; X_Im[136]=-32'd0; X_Im[137]=-32'd0; X_Im[138]=-32'd0; X_Im[139]=-32'd0; X_Im[140]=-32'd0; X_Im[141]=-32'd0; X_Im[142]=-32'd0; X_Im[143]=-32'd0; X_Im[144]=32'd0; X_Im[145]=32'd0; X_Im[146]=32'd0; X_Im[147]=32'd0; X_Im[148]=32'd0; X_Im[149]=32'd0; X_Im[150]=32'd0; X_Im[151]=-32'd0; X_Im[152]=32'd0; X_Im[153]=32'd0; X_Im[154]=32'd0; X_Im[155]=-32'd0; X_Im[156]=-32'd0; X_Im[157]=-32'd0; X_Im[158]=32'd0; X_Im[159]=32'd0; X_Im[160]=32'd0; X_Im[161]=32'd0; X_Im[162]=32'd0; X_Im[163]=-32'd0; X_Im[164]=-32'd0; X_Im[165]=-32'd0; X_Im[166]=-32'd0; X_Im[167]=-32'd0; X_Im[168]=-32'd0; X_Im[169]=-32'd0; X_Im[170]=-32'd0; X_Im[171]=32'd0; X_Im[172]=-32'd0; X_Im[173]=32'd0; X_Im[174]=32'd0; X_Im[175]=32'd0; X_Im[176]=32'd0; X_Im[177]=32'd0; X_Im[178]=32'd0; X_Im[179]=32'd0; X_Im[180]=32'd0; X_Im[181]=-32'd0; X_Im[182]=-32'd0; X_Im[183]=-32'd0; X_Im[184]=32'd0; X_Im[185]=32'd0; X_Im[186]=32'd0; X_Im[187]=32'd0; X_Im[188]=-32'd0; X_Im[189]=-32'd0; X_Im[190]=-32'd0; X_Im[191]=-32'd0; X_Im[192]=-32'd0; X_Im[193]=32'd0; X_Im[194]=32'd0; X_Im[195]=32'd0; X_Im[196]=-32'd0; X_Im[197]=-32'd0; X_Im[198]=-32'd0; X_Im[199]=32'd0; X_Im[200]=32'd0; X_Im[201]=32'd0; X_Im[202]=32'd0; X_Im[203]=32'd0; X_Im[204]=32'd0; X_Im[205]=32'd0; X_Im[206]=32'd0; X_Im[207]=32'd0; X_Im[208]=32'd0; X_Im[209]=32'd0; X_Im[210]=32'd0; X_Im[211]=32'd0; X_Im[212]=32'd0; X_Im[213]=-32'd0; X_Im[214]=-32'd0; X_Im[215]=-32'd0; X_Im[216]=-32'd0; X_Im[217]=-32'd0; X_Im[218]=-32'd0; X_Im[219]=-32'd0; X_Im[220]=-32'd0; X_Im[221]=-32'd0; X_Im[222]=-32'd0; X_Im[223]=-32'd0; X_Im[224]=-32'd0; X_Im[225]=-32'd0; X_Im[226]=32'd0; X_Im[227]=32'd0; X_Im[228]=32'd0; X_Im[229]=32'd0; X_Im[230]=32'd0; X_Im[231]=32'd0; X_Im[232]=32'd0; X_Im[233]=32'd0; X_Im[234]=-32'd0; X_Im[235]=-32'd0; X_Im[236]=32'd0; X_Im[237]=32'd0; X_Im[238]=32'd0; X_Im[239]=32'd0; X_Im[240]=-32'd0; X_Im[241]=-32'd0; X_Im[242]=-32'd0; X_Im[243]=-32'd0; X_Im[244]=-32'd0; X_Im[245]=-32'd0; X_Im[246]=-32'd0; X_Im[247]=32'd0; X_Im[248]=32'd0; X_Im[249]=32'd0; X_Im[250]=32'd0; X_Im[251]=32'd0; X_Im[252]=32'd0; X_Im[253]=32'd0; X_Im[254]=32'd0; X_Im[255]=32'd0; X_Im[256]=32'd0; X_Im[257]=-32'd0; X_Im[258]=-32'd0; X_Im[259]=-32'd0; X_Im[260]=32'd0; X_Im[261]=32'd0; X_Im[262]=32'd0; X_Im[263]=32'd0; X_Im[264]=32'd0; X_Im[265]=32'd0; X_Im[266]=32'd0; X_Im[267]=-32'd0; X_Im[268]=-32'd0; X_Im[269]=-32'd0; X_Im[270]=-32'd0; X_Im[271]=-32'd0; X_Im[272]=-32'd0; X_Im[273]=-32'd0; X_Im[274]=-32'd0; X_Im[275]=-32'd0; X_Im[276]=32'd0; X_Im[277]=32'd0; X_Im[278]=32'd0; X_Im[279]=32'd0; X_Im[280]=32'd0; X_Im[281]=32'd0; X_Im[282]=32'd0; X_Im[283]=32'd0; X_Im[284]=32'd0; X_Im[285]=32'd0; X_Im[286]=32'd0; X_Im[287]=32'd0; X_Im[288]=32'd0; X_Im[289]=-32'd0; X_Im[290]=-32'd0; X_Im[291]=-32'd0; X_Im[292]=-32'd0; X_Im[293]=32'd0; X_Im[294]=-32'd0; X_Im[295]=-32'd0; X_Im[296]=-32'd0; X_Im[297]=-32'd0; X_Im[298]=-32'd0; X_Im[299]=32'd0; X_Im[300]=32'd0; X_Im[301]=32'd0; X_Im[302]=-32'd0; X_Im[303]=-32'd0; X_Im[304]=-32'd0; X_Im[305]=-32'd0; X_Im[306]=32'd0; X_Im[307]=32'd0; X_Im[308]=32'd0; X_Im[309]=32'd0; X_Im[310]=32'd0; X_Im[311]=-32'd0; X_Im[312]=32'd0; X_Im[313]=32'd0; X_Im[314]=32'd0; X_Im[315]=32'd0; X_Im[316]=32'd0; X_Im[317]=-32'd0; X_Im[318]=-32'd0; X_Im[319]=-32'd0; X_Im[320]=-32'd0; X_Im[321]=-32'd0; X_Im[322]=-32'd0; X_Im[323]=-32'd0; X_Im[324]=-32'd0; X_Im[325]=-32'd0; X_Im[326]=-32'd0; X_Im[327]=-32'd0; X_Im[328]=-32'd0; X_Im[329]=32'd0; X_Im[330]=32'd0; X_Im[331]=32'd0; X_Im[332]=32'd0; X_Im[333]=32'd0; X_Im[334]=32'd0; X_Im[335]=-32'd0; X_Im[336]=-32'd0; X_Im[337]=-32'd0; X_Im[338]=32'd0; X_Im[339]=32'd0; X_Im[340]=32'd0; X_Im[341]=32'd0; X_Im[342]=-32'd0; X_Im[343]=-32'd0; X_Im[344]=-32'd0; X_Im[345]=-32'd0; X_Im[346]=-32'd0; X_Im[347]=-32'd0; X_Im[348]=-32'd0; X_Im[349]=-32'd0; X_Im[350]=-32'd0; X_Im[351]=-32'd0; X_Im[352]=32'd0; X_Im[353]=32'd0; X_Im[354]=32'd0; X_Im[355]=32'd0; X_Im[356]=32'd0; X_Im[357]=32'd0; X_Im[358]=32'd0; X_Im[359]=32'd0; X_Im[360]=32'd0; X_Im[361]=32'd0; X_Im[362]=32'd0; X_Im[363]=32'd0; X_Im[364]=32'd0; X_Im[365]=32'd0; X_Im[366]=32'd0; X_Im[367]=32'd0; X_Im[368]=32'd0; X_Im[369]=32'd0; X_Im[370]=32'd0; X_Im[371]=-32'd0; X_Im[372]=-32'd0; X_Im[373]=-32'd0; X_Im[374]=-32'd0; X_Im[375]=-32'd0; X_Im[376]=-32'd0; X_Im[377]=-32'd0; X_Im[378]=-32'd0; X_Im[379]=-32'd0; X_Im[380]=-32'd0; X_Im[381]=-32'd0; X_Im[382]=32'd0; X_Im[383]=32'd0; X_Im[384]=32'd0; X_Im[385]=32'd0; X_Im[386]=32'd0; X_Im[387]=32'd0; X_Im[388]=32'd0; X_Im[389]=32'd0; X_Im[390]=32'd0; X_Im[391]=32'd0; X_Im[392]=32'd0; X_Im[393]=-32'd0; X_Im[394]=-32'd0; X_Im[395]=-32'd0; X_Im[396]=-32'd0; X_Im[397]=-32'd0; X_Im[398]=-32'd0; X_Im[399]=32'd0; X_Im[400]=32'd0; X_Im[401]=32'd0; X_Im[402]=32'd0; X_Im[403]=32'd0; X_Im[404]=32'd0; X_Im[405]=32'd0; X_Im[406]=32'd0; X_Im[407]=32'd0; X_Im[408]=32'd0; X_Im[409]=32'd0; X_Im[410]=32'd0; X_Im[411]=-32'd0; X_Im[412]=-32'd0; X_Im[413]=32'd0; X_Im[414]=32'd0; X_Im[415]=32'd0; X_Im[416]=32'd0; X_Im[417]=32'd0; X_Im[418]=32'd0; X_Im[419]=32'd0; X_Im[420]=-32'd0; X_Im[421]=-32'd0; X_Im[422]=-32'd0; X_Im[423]=-32'd0; X_Im[424]=-32'd0; X_Im[425]=-32'd0; X_Im[426]=-32'd0; X_Im[427]=-32'd0; X_Im[428]=-32'd0; X_Im[429]=-32'd0; X_Im[430]=32'd0; X_Im[431]=32'd0; X_Im[432]=32'd0; X_Im[433]=32'd0; X_Im[434]=32'd0; X_Im[435]=32'd0; X_Im[436]=32'd0; X_Im[437]=32'd0; X_Im[438]=32'd0; X_Im[439]=32'd0; X_Im[440]=-32'd0; X_Im[441]=-32'd0; X_Im[442]=-32'd0; X_Im[443]=32'd0; X_Im[444]=32'd0; X_Im[445]=32'd0; X_Im[446]=32'd0; X_Im[447]=32'd0; X_Im[448]=32'd0; X_Im[449]=-32'd0; X_Im[450]=-32'd0; X_Im[451]=-32'd0; X_Im[452]=-32'd0; X_Im[453]=-32'd0; X_Im[454]=-32'd0; X_Im[455]=-32'd0; X_Im[456]=-32'd0; X_Im[457]=-32'd0; X_Im[458]=-32'd0; X_Im[459]=32'd0; X_Im[460]=32'd0; X_Im[461]=32'd0; X_Im[462]=32'd0; X_Im[463]=32'd0; X_Im[464]=32'd0; X_Im[465]=32'd0; X_Im[466]=-32'd0; X_Im[467]=32'd0; X_Im[468]=32'd0; X_Im[469]=32'd0; X_Im[470]=-32'd0; X_Im[471]=-32'd0; X_Im[472]=-32'd0; X_Im[473]=-32'd0; X_Im[474]=-32'd0; X_Im[475]=-32'd0; X_Im[476]=-32'd0; X_Im[477]=-32'd0; X_Im[478]=-32'd0; X_Im[479]=-32'd0; X_Im[480]=-32'd0; X_Im[481]=-32'd0; X_Im[482]=-32'd0; X_Im[483]=-32'd0; X_Im[484]=-32'd0; X_Im[485]=-32'd0; X_Im[486]=32'd0; X_Im[487]=32'd0; X_Im[488]=-32'd0; X_Im[489]=32'd0; X_Im[490]=32'd0; X_Im[491]=32'd0; X_Im[492]=32'd0; X_Im[493]=32'd0; X_Im[494]=32'd0; X_Im[495]=32'd0; X_Im[496]=-32'd0; X_Im[497]=-32'd0; X_Im[498]=-32'd0; X_Im[499]=-32'd0; X_Im[500]=-32'd0; X_Im[501]=-32'd0; X_Im[502]=-32'd0; X_Im[503]=-32'd0; X_Im[504]=-32'd0; X_Im[505]=-32'd0; X_Im[506]=32'd0; X_Im[507]=32'd0; X_Im[508]=32'd0; X_Im[509]=32'd0; X_Im[510]=32'd0; X_Im[511]=32'd0; X_Im[512]=32'd0; X_Im[513]=-32'd0; X_Im[514]=-32'd0; X_Im[515]=32'd0; X_Im[516]=-32'd0; X_Im[517]=32'd0; X_Im[518]=32'd0; X_Im[519]=32'd0; X_Im[520]=32'd0; X_Im[521]=32'd0; X_Im[522]=32'd0; X_Im[523]=32'd0; X_Im[524]=32'd0; X_Im[525]=32'd0; X_Im[526]=-32'd0; X_Im[527]=-32'd0; X_Im[528]=-32'd0; X_Im[529]=-32'd0; X_Im[530]=-32'd0; X_Im[531]=-32'd0; X_Im[532]=-32'd0; X_Im[533]=-32'd0; X_Im[534]=-32'd0; X_Im[535]=32'd0; X_Im[536]=32'd0; X_Im[537]=32'd0; X_Im[538]=32'd0; X_Im[539]=32'd0; X_Im[540]=32'd0; X_Im[541]=32'd0; X_Im[542]=32'd0; X_Im[543]=32'd0; X_Im[544]=32'd0; X_Im[545]=32'd0; X_Im[546]=-32'd0; X_Im[547]=-32'd0; X_Im[548]=-32'd0; X_Im[549]=-32'd0; X_Im[550]=-32'd0; X_Im[551]=32'd0; X_Im[552]=32'd0; X_Im[553]=32'd0; X_Im[554]=32'd0; X_Im[555]=32'd0; X_Im[556]=32'd0; X_Im[557]=32'd0; X_Im[558]=-32'd0; X_Im[559]=-32'd0; X_Im[560]=-32'd0; X_Im[561]=-32'd0; X_Im[562]=-32'd0; X_Im[563]=-32'd0; X_Im[564]=-32'd0; X_Im[565]=-32'd0; X_Im[566]=32'd0; X_Im[567]=32'd0; X_Im[568]=32'd0; X_Im[569]=32'd0; X_Im[570]=32'd0; X_Im[571]=32'd0; X_Im[572]=32'd0; X_Im[573]=-32'd0; X_Im[574]=-32'd0; X_Im[575]=-32'd0; X_Im[576]=-32'd0; X_Im[577]=-32'd0; X_Im[578]=-32'd0; X_Im[579]=-32'd0; X_Im[580]=-32'd0; X_Im[581]=-32'd0; X_Im[582]=-32'd0; X_Im[583]=-32'd0; X_Im[584]=-32'd0; X_Im[585]=32'd0; X_Im[586]=32'd0; X_Im[587]=32'd0; X_Im[588]=32'd0; X_Im[589]=32'd0; X_Im[590]=32'd0; X_Im[591]=32'd0; X_Im[592]=-32'd0; X_Im[593]=-32'd0; X_Im[594]=-32'd0; X_Im[595]=-32'd0; X_Im[596]=32'd0; X_Im[597]=32'd0; X_Im[598]=32'd0; X_Im[599]=32'd0; X_Im[600]=32'd0; X_Im[601]=32'd0; X_Im[602]=32'd0; X_Im[603]=32'd0; X_Im[604]=-32'd0; X_Im[605]=-32'd0; X_Im[606]=-32'd0; X_Im[607]=-32'd0; X_Im[608]=-32'd0; X_Im[609]=-32'd0; X_Im[610]=-32'd0; X_Im[611]=-32'd0; X_Im[612]=-32'd0; X_Im[613]=32'd0; X_Im[614]=32'd0; X_Im[615]=32'd0; X_Im[616]=32'd0; X_Im[617]=32'd0; X_Im[618]=32'd0; X_Im[619]=32'd0; X_Im[620]=32'd0; X_Im[621]=32'd0; X_Im[622]=-32'd0; X_Im[623]=-32'd0; X_Im[624]=32'd0; X_Im[625]=-32'd0; X_Im[626]=-32'd0; X_Im[627]=32'd0; X_Im[628]=32'd0; X_Im[629]=32'd0; X_Im[630]=32'd0; X_Im[631]=-32'd0; X_Im[632]=-32'd0; X_Im[633]=-32'd0; X_Im[634]=-32'd0; X_Im[635]=-32'd0; X_Im[636]=-32'd0; X_Im[637]=-32'd0; X_Im[638]=-32'd0; X_Im[639]=-32'd0; X_Im[640]=32'd0; X_Im[641]=32'd0; X_Im[642]=32'd0; X_Im[643]=32'd0; X_Im[644]=32'd0; X_Im[645]=32'd0; X_Im[646]=32'd0; X_Im[647]=32'd0; X_Im[648]=32'd0; X_Im[649]=32'd0; X_Im[650]=32'd0; X_Im[651]=-32'd0; X_Im[652]=-32'd0; X_Im[653]=-32'd0; X_Im[654]=-32'd0; X_Im[655]=-32'd0; X_Im[656]=-32'd0; X_Im[657]=-32'd0; X_Im[658]=-32'd0; X_Im[659]=32'd0; X_Im[660]=32'd0; X_Im[661]=32'd0; X_Im[662]=32'd0; X_Im[663]=32'd0; X_Im[664]=32'd0; X_Im[665]=32'd0; X_Im[666]=-32'd0; X_Im[667]=-32'd0; X_Im[668]=-32'd0; X_Im[669]=-32'd0; X_Im[670]=-32'd0; X_Im[671]=32'd0; X_Im[672]=32'd0; X_Im[673]=32'd0; X_Im[674]=32'd0; X_Im[675]=32'd0; X_Im[676]=32'd0; X_Im[677]=32'd0; X_Im[678]=32'd0; X_Im[679]=32'd0; X_Im[680]=32'd0; X_Im[681]=-32'd0; X_Im[682]=-32'd0; X_Im[683]=-32'd0; X_Im[684]=-32'd0; X_Im[685]=-32'd0; X_Im[686]=-32'd0; X_Im[687]=-32'd0; X_Im[688]=-32'd0; X_Im[689]=-32'd0; X_Im[690]=32'd0; X_Im[691]=32'd0; X_Im[692]=32'd0; X_Im[693]=32'd0; X_Im[694]=32'd0; X_Im[695]=32'd0; X_Im[696]=32'd0; X_Im[697]=-32'd0; X_Im[698]=-32'd0; X_Im[699]=-32'd0; X_Im[700]=-32'd0; X_Im[701]=-32'd0; X_Im[702]=-32'd0; X_Im[703]=-32'd0; X_Im[704]=-32'd0; X_Im[705]=32'd0; X_Im[706]=32'd0; X_Im[707]=32'd0; X_Im[708]=32'd0; X_Im[709]=32'd0; X_Im[710]=32'd0; X_Im[711]=-32'd0; X_Im[712]=-32'd0; X_Im[713]=-32'd0; X_Im[714]=-32'd0; X_Im[715]=-32'd0; X_Im[716]=-32'd0; X_Im[717]=-32'd0; X_Im[718]=-32'd0; X_Im[719]=32'd0; X_Im[720]=32'd0; X_Im[721]=32'd0; X_Im[722]=32'd0; X_Im[723]=32'd0; X_Im[724]=32'd0; X_Im[725]=32'd0; X_Im[726]=32'd0; X_Im[727]=32'd0; X_Im[728]=-32'd0; X_Im[729]=-32'd0; X_Im[730]=-32'd0; X_Im[731]=-32'd0; X_Im[732]=-32'd0; X_Im[733]=-32'd0; X_Im[734]=-32'd0; X_Im[735]=-32'd0; X_Im[736]=-32'd0; X_Im[737]=-32'd0; X_Im[738]=-32'd0; X_Im[739]=32'd0; X_Im[740]=32'd0; X_Im[741]=32'd0; X_Im[742]=-32'd0; X_Im[743]=-32'd0; X_Im[744]=32'd0; X_Im[745]=32'd0; X_Im[746]=32'd0; X_Im[747]=32'd0; X_Im[748]=32'd0; X_Im[749]=32'd0; X_Im[750]=32'd0; X_Im[751]=32'd0; X_Im[752]=32'd0; X_Im[753]=32'd0; X_Im[754]=32'd0; X_Im[755]=32'd0; X_Im[756]=32'd0; X_Im[757]=32'd0; X_Im[758]=-32'd0; X_Im[759]=-32'd0; X_Im[760]=-32'd0; X_Im[761]=-32'd0; X_Im[762]=-32'd0; X_Im[763]=-32'd0; X_Im[764]=-32'd0; X_Im[765]=32'd0; X_Im[766]=32'd0; X_Im[767]=32'd0; X_Im[768]=32'd0; X_Im[769]=32'd0; X_Im[770]=32'd0; X_Im[771]=32'd0; X_Im[772]=32'd0; X_Im[773]=32'd0; X_Im[774]=-32'd0; X_Im[775]=-32'd0; X_Im[776]=-32'd0; X_Im[777]=-32'd0; X_Im[778]=-32'd0; X_Im[779]=32'd0; X_Im[780]=32'd0; X_Im[781]=32'd0; X_Im[782]=32'd0; X_Im[783]=32'd0; X_Im[784]=32'd0; X_Im[785]=32'd0; X_Im[786]=32'd0; X_Im[787]=-32'd0; X_Im[788]=-32'd0; X_Im[789]=-32'd0; X_Im[790]=-32'd0; X_Im[791]=-32'd0; X_Im[792]=-32'd0; X_Im[793]=-32'd0; X_Im[794]=-32'd0; X_Im[795]=32'd0; X_Im[796]=32'd0; X_Im[797]=32'd0; X_Im[798]=32'd0; X_Im[799]=32'd0; X_Im[800]=32'd0; X_Im[801]=32'd0; X_Im[802]=32'd0; X_Im[803]=-32'd0; X_Im[804]=-32'd0; X_Im[805]=-32'd0; X_Im[806]=-32'd0; X_Im[807]=-32'd0; X_Im[808]=-32'd0; X_Im[809]=-32'd0; X_Im[810]=32'd0; X_Im[811]=32'd0; X_Im[812]=-32'd0; X_Im[813]=32'd0; X_Im[814]=32'd0; X_Im[815]=32'd0; X_Im[816]=32'd0; X_Im[817]=32'd0; X_Im[818]=-32'd0; X_Im[819]=-32'd0; X_Im[820]=-32'd0; X_Im[821]=-32'd0; X_Im[822]=-32'd0; X_Im[823]=-32'd0; X_Im[824]=32'd0; X_Im[825]=32'd0; X_Im[826]=32'd0; X_Im[827]=32'd0; X_Im[828]=32'd0; X_Im[829]=32'd0; X_Im[830]=32'd0; X_Im[831]=32'd0; X_Im[832]=32'd0; X_Im[833]=32'd0; X_Im[834]=32'd0; X_Im[835]=-32'd0; X_Im[836]=-32'd0; X_Im[837]=-32'd0; X_Im[838]=-32'd0; X_Im[839]=-32'd0; X_Im[840]=-32'd0; X_Im[841]=-32'd0; X_Im[842]=32'd0; X_Im[843]=32'd0; X_Im[844]=32'd0; X_Im[845]=32'd0; X_Im[846]=32'd0; X_Im[847]=32'd0; X_Im[848]=32'd0; X_Im[849]=32'd0; X_Im[850]=32'd0; X_Im[851]=-32'd0; X_Im[852]=-32'd0; X_Im[853]=-32'd0; X_Im[854]=-32'd0; X_Im[855]=-32'd0; X_Im[856]=32'd0; X_Im[857]=32'd0; X_Im[858]=32'd0; X_Im[859]=32'd0; X_Im[860]=32'd0; X_Im[861]=32'd0; X_Im[862]=32'd0; X_Im[863]=32'd0; X_Im[864]=-32'd0; X_Im[865]=-32'd0; X_Im[866]=-32'd0; X_Im[867]=-32'd0; X_Im[868]=-32'd0; X_Im[869]=-32'd0; X_Im[870]=-32'd0; X_Im[871]=-32'd0; X_Im[872]=-32'd0; X_Im[873]=-32'd0; X_Im[874]=32'd0; X_Im[875]=32'd0; X_Im[876]=32'd0; X_Im[877]=32'd0; X_Im[878]=32'd0; X_Im[879]=32'd0; X_Im[880]=-32'd0; X_Im[881]=-32'd0; X_Im[882]=-32'd0; X_Im[883]=-32'd0; X_Im[884]=32'd0; X_Im[885]=32'd0; X_Im[886]=32'd0; X_Im[887]=32'd0; X_Im[888]=32'd0; X_Im[889]=-32'd0; X_Im[890]=-32'd0; X_Im[891]=-32'd0; X_Im[892]=32'd0; X_Im[893]=32'd0; X_Im[894]=32'd0; X_Im[895]=-32'd0; X_Im[896]=-32'd0; X_Im[897]=-32'd0; X_Im[898]=-32'd0; X_Im[899]=-32'd0; X_Im[900]=32'd0; X_Im[901]=32'd0; X_Im[902]=32'd0; X_Im[903]=32'd0; X_Im[904]=32'd0; X_Im[905]=32'd0; X_Im[906]=32'd0; X_Im[907]=32'd0; X_Im[908]=32'd0; X_Im[909]=32'd0; X_Im[910]=32'd0; X_Im[911]=-32'd0; X_Im[912]=-32'd0; X_Im[913]=-32'd0; X_Im[914]=-32'd0; X_Im[915]=-32'd0; X_Im[916]=-32'd0; X_Im[917]=-32'd0; X_Im[918]=-32'd0; X_Im[919]=-32'd0; X_Im[920]=-32'd0; X_Im[921]=-32'd0; X_Im[922]=-32'd0; X_Im[923]=32'd0; X_Im[924]=32'd0; X_Im[925]=32'd0; X_Im[926]=32'd0; X_Im[927]=32'd0; X_Im[928]=-32'd0; X_Im[929]=-32'd0; X_Im[930]=-32'd0; X_Im[931]=-32'd0; X_Im[932]=-32'd0; X_Im[933]=-32'd0; X_Im[934]=32'd0; X_Im[935]=32'd0; X_Im[936]=32'd0; X_Im[937]=32'd0; X_Im[938]=32'd0; X_Im[939]=32'd0; X_Im[940]=32'd0; X_Im[941]=-32'd0; X_Im[942]=-32'd0; X_Im[943]=-32'd0; X_Im[944]=-32'd0; X_Im[945]=-32'd0; X_Im[946]=-32'd0; X_Im[947]=-32'd0; X_Im[948]=-32'd0; X_Im[949]=32'd0; X_Im[950]=32'd0; X_Im[951]=32'd0; X_Im[952]=32'd0; X_Im[953]=32'd0; X_Im[954]=32'd0; X_Im[955]=32'd0; X_Im[956]=32'd0; X_Im[957]=-32'd0; X_Im[958]=-32'd0; X_Im[959]=-32'd0; X_Im[960]=-32'd0; X_Im[961]=-32'd0; X_Im[962]=-32'd0; X_Im[963]=32'd0; X_Im[964]=32'd0; X_Im[965]=32'd0; X_Im[966]=32'd0; X_Im[967]=32'd0; X_Im[968]=32'd0; X_Im[969]=32'd0; X_Im[970]=32'd0; X_Im[971]=32'd0; X_Im[972]=-32'd0; X_Im[973]=-32'd0; X_Im[974]=-32'd0; X_Im[975]=-32'd0; X_Im[976]=-32'd0; X_Im[977]=-32'd0; X_Im[978]=-32'd0; X_Im[979]=32'd0; X_Im[980]=32'd0; X_Im[981]=32'd0; X_Im[982]=32'd0; X_Im[983]=32'd0; X_Im[984]=32'd0; X_Im[985]=32'd0; X_Im[986]=32'd0; X_Im[987]=32'd0; X_Im[988]=-32'd0; X_Im[989]=-32'd0; X_Im[990]=-32'd0; X_Im[991]=-32'd0; X_Im[992]=-32'd0; X_Im[993]=-32'd0; X_Im[994]=-32'd0; X_Im[995]=-32'd0; X_Im[996]=32'd0; X_Im[997]=32'd0; X_Im[998]=32'd0; X_Im[999]=32'd0; X_Im[1000]=32'd0; X_Im[1001]=32'd0; X_Im[1002]=32'd0; X_Im[1003]=-32'd0; X_Im[1004]=-32'd0; X_Im[1005]=-32'd0; X_Im[1006]=-32'd0; X_Im[1007]=-32'd0; X_Im[1008]=-32'd0; X_Im[1009]=-32'd0; X_Im[1010]=-32'd0; X_Im[1011]=32'd0; X_Im[1012]=32'd0; X_Im[1013]=32'd0; X_Im[1014]=32'd0; X_Im[1015]=32'd0; X_Im[1016]=32'd0; X_Im[1017]=32'd0; X_Im[1018]=32'd0; X_Im[1019]=-32'd0; X_Im[1020]=-32'd0; X_Im[1021]=-32'd0; X_Im[1022]=-32'd0; X_Im[1023]=-32'd0;
		#10
		Reset = 0;
		#10
		
		Start = 1;
		#130
		Start = 0;
	end

endmodule