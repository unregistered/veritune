`timescale 1ns / 1ps

module IFFT1024_tb_v;
	parameter PRE = 32;
		
	reg Clk;
	reg Reset, Start, Ack;
	reg signed [PRE-1:0] X_Re [1023:0];
	reg signed [PRE-1:0] X_Im [1023:0];
	integer timestamp;
	
	// Outputs
	wire [3:0] state;
	wire Done;
	wire signed [31:0] x_top_re;
	wire signed [31:0] x_top_im;
	wire signed [31:0] x_bot_re;
	wire signed [31:0] x_bot_im;	
	wire signed [31:0] x_re_0, x_re_1, x_re_2, x_re_3, x_re_4, x_re_5, x_re_6, x_re_7;
	wire signed [31:0] x_im_0, x_im_1, x_im_2, x_im_3, x_im_4, x_im_5, x_im_6, x_im_7;
	assign x_re_0 = X_Re[0];
	assign x_re_1 = X_Re[1];
	assign x_re_2 = X_Re[2];
	assign x_re_3 = X_Re[3];
	assign x_re_4 = X_Re[4];
	assign x_re_5 = X_Re[5];
	assign x_re_6 = X_Re[6];
	assign x_re_7 = X_Re[7];
	assign x_im_0 = X_Im[0];
	assign x_im_1 = X_Im[1];
	assign x_im_2 = X_Im[2];
	assign x_im_3 = X_Im[3];
	assign x_im_4 = X_Im[4];
	assign x_im_5 = X_Im[5];
	assign x_im_6 = X_Im[6];
	assign x_im_7 = X_Im[7];	
	
	// Internal
	wire signed [31:0] y_top_re;
	wire signed [31:0] y_top_im;
	wire signed [31:0] y_bot_re;
	wire signed [31:0] y_bot_im;
	wire [9:0]  i_top, i_bot;
	assign x_top_re = X_Re[i_top];
	assign x_top_im = X_Im[i_top];
	assign x_bot_re = X_Re[i_bot];
	assign x_bot_im = X_Im[i_bot];
	
		
	
	// Instantiate the Unit Under Test (UUT)
	FFT1024 uut_ifft (
		//	Ins
		.Clk(Clk),
		.Reset(Reset),
		.Start(Start),
		.Ack(Ack),
		// Swap the reals and ims
		.x_top_re(X_Im[i_top]),
		.x_top_im(X_Re[i_top]),
		.x_bot_re(X_Im[i_bot]),
		.x_bot_im(X_Re[i_bot]),
		//	Outs
		.i_top(i_top),
		.i_bot(i_bot),
		// Swap reals and ims
		.y_top_re(y_top_im),
		.y_top_im(y_top_re),
		.y_bot_re(y_bot_im),
		.y_bot_im(y_bot_re),
		.Done(Done),
		.state(state)
	);
	
	
	initial
	begin
		Clk = 0; // Initialize clock
		Start = 0;
		Reset = 0;
	end
	
	// Keep clock running
	always
	begin
		#20; 
		Clk = ~ Clk; 
	end
	
	//	Here's how to use the butterfly unit
	always @(posedge Clk)
	begin
		timestamp <= timestamp + 1;
		case(state)
			4'd1: //Done
			begin
				$display("X[0]=%d + i%d", X_Re[0]>>>10, X_Im[0]>>>10);
				$display("X[1]=%d + i%d", X_Re[1]>>>10, X_Im[1]>>>10);
				$display("X[2]=%d + i%d", X_Re[2]>>>10, X_Im[2]>>>10);
				$display("X[3]=%d + i%d", X_Re[3]>>>10, X_Im[3]>>>10);
				$display("X[4]=%d + i%d", X_Re[4]>>>10, X_Im[4]>>>10);
				$display("X[5]=%d + i%d", X_Re[5]>>>10, X_Im[5]>>>10);
				$display("X[6]=%d + i%d", X_Re[6]>>>10, X_Im[6]>>>10);
				$display("X[7]=%d + i%d", X_Re[7]>>>10, X_Im[7]>>>10);
				Ack = 1;
			end
			4'd2: //Proc
			begin
				$display("Time: %d", timestamp);
				$display("  i_top %b i_bot %b", i_top, i_bot);
				$display("  x_top_re %d x_bot_re %d", X_Re[i_top], X_Re[i_bot]);
				$display("  y_top %d + i%d y_bot %d + i%d", y_top_re, y_top_im, y_bot_re, y_bot_im);
				X_Re[i_top] <= y_top_re;
				X_Im[i_top] <= y_top_im;
				X_Re[i_bot] <= y_bot_re;
				X_Im[i_bot] <= y_bot_im;
			end
		endcase
	end
	
	//	Just setup
	initial
	begin
		timestamp = 0;
		Start = 0;
		Reset = 0;
		Ack = 0;
		#10
		Reset = 1;
		#200
		// IFFT
		X_Re[0]=32'd87845; X_Re[512]=32'd3344; X_Re[256]=32'd8055; X_Re[768]=-32'd3237; X_Re[128]=-32'd3178; X_Re[640]=-32'd8097; X_Re[384]=-32'd13493; X_Re[896]=-32'd45742; X_Re[64]=-32'd5662; X_Re[576]=-32'd166613; X_Re[320]=-32'd45666; X_Re[832]=32'd71943; X_Re[192]=-32'd7187; X_Re[704]=-32'd40016; X_Re[448]=32'd2080; X_Re[960]=32'd16013; X_Re[32]=-32'd12426; X_Re[544]=32'd41019; X_Re[288]=-32'd32079; X_Re[800]=-32'd54871; X_Re[160]=32'd1037; X_Re[672]=-32'd19342; X_Re[416]=-32'd4748; X_Re[928]=32'd13800; X_Re[96]=-32'd5577; X_Re[608]=32'd2592; X_Re[352]=32'd41646; X_Re[864]=-32'd73347; X_Re[224]=-32'd34797; X_Re[736]=-32'd23890; X_Re[480]=-32'd38433; X_Re[992]=-32'd23713; X_Re[16]=-32'd20014; X_Re[528]=-32'd10798; X_Re[272]=-32'd22086; X_Re[784]=32'd31774; X_Re[144]=-32'd57943; X_Re[656]=-32'd33674; X_Re[400]=-32'd92155; X_Re[912]=-32'd219111; X_Re[80]=32'd422815; X_Re[592]=32'd77266; X_Re[336]=32'd48085; X_Re[848]=32'd19080; X_Re[208]=32'd71278; X_Re[720]=32'd32371; X_Re[464]=32'd7926; X_Re[976]=32'd35091; X_Re[48]=32'd37484; X_Re[560]=32'd19509; X_Re[304]=32'd18707; X_Re[816]=32'd44296; X_Re[176]=32'd3041; X_Re[688]=32'd200812; X_Re[432]=-32'd32042; X_Re[944]=-32'd2465; X_Re[112]=32'd19028; X_Re[624]=32'd16164; X_Re[368]=32'd99801; X_Re[880]=32'd172680; X_Re[240]=-32'd374488; X_Re[752]=-32'd76563; X_Re[496]=-32'd68355; X_Re[1008]=-32'd73725; X_Re[8]=-32'd89550; X_Re[520]=-32'd84078; X_Re[264]=-32'd350559; X_Re[776]=-32'd220475; X_Re[136]=32'd25897; X_Re[648]=32'd98286; X_Re[392]=32'd24689; X_Re[904]=32'd86424; X_Re[72]=32'd20529; X_Re[584]=32'd27560; X_Re[328]=32'd24094; X_Re[840]=32'd20953; X_Re[200]=32'd15514; X_Re[712]=32'd18835; X_Re[456]=-32'd2159; X_Re[968]=-32'd322659; X_Re[40]=-32'd103143; X_Re[552]=32'd21865; X_Re[296]=32'd5014; X_Re[808]=32'd10478; X_Re[168]=32'd7487; X_Re[680]=32'd1599; X_Re[424]=32'd508; X_Re[936]=32'd6553; X_Re[104]=32'd12647; X_Re[616]=32'd328; X_Re[360]=32'd13322; X_Re[872]=32'd19519; X_Re[232]=32'd10361; X_Re[744]=32'd11635; X_Re[488]=32'd53368; X_Re[1000]=-32'd32083; X_Re[24]=-32'd1423; X_Re[536]=-32'd15483; X_Re[280]=-32'd6194; X_Re[792]=32'd3784; X_Re[152]=32'd2743; X_Re[664]=32'd2850; X_Re[408]=-32'd429; X_Re[920]=-32'd6999; X_Re[88]=-32'd8783; X_Re[600]=-32'd33732; X_Re[344]=32'd36890; X_Re[856]=32'd20766; X_Re[216]=32'd2968; X_Re[728]=32'd13462; X_Re[472]=-32'd870; X_Re[984]=32'd7264; X_Re[56]=-32'd4449; X_Re[568]=32'd4331; X_Re[312]=32'd8206; X_Re[824]=32'd3472; X_Re[184]=32'd7848; X_Re[696]=32'd24008; X_Re[440]=-32'd14034; X_Re[952]=-32'd93185; X_Re[120]=32'd35868; X_Re[632]=-32'd8956; X_Re[376]=32'd16199; X_Re[888]=32'd4346; X_Re[248]=-32'd653; X_Re[760]=32'd11710; X_Re[504]=32'd242; X_Re[1016]=-32'd2025; X_Re[4]=-32'd2026; X_Re[516]=-32'd5956; X_Re[260]=32'd1626; X_Re[772]=-32'd5217; X_Re[132]=32'd28921; X_Re[644]=32'd348596; X_Re[388]=32'd70108; X_Re[900]=-32'd59599; X_Re[68]=32'd4423; X_Re[580]=-32'd10221; X_Re[324]=-32'd2938; X_Re[836]=-32'd7719; X_Re[196]=-32'd14770; X_Re[708]=32'd24684; X_Re[452]=32'd8862; X_Re[964]=-32'd7572; X_Re[36]=32'd2346; X_Re[548]=32'd1621; X_Re[292]=32'd7001; X_Re[804]=32'd5648; X_Re[164]=32'd1191; X_Re[676]=32'd3541; X_Re[420]=32'd8099; X_Re[932]=32'd9251; X_Re[100]=32'd4481; X_Re[612]=32'd5927; X_Re[356]=-32'd785; X_Re[868]=32'd7908; X_Re[228]=-32'd9583; X_Re[740]=32'd16551; X_Re[484]=32'd43192; X_Re[996]=-32'd26098; X_Re[20]=32'd44207; X_Re[532]=-32'd53731; X_Re[276]=-32'd13945; X_Re[788]=32'd7595; X_Re[148]=-32'd18047; X_Re[660]=-32'd7142; X_Re[404]=32'd2843; X_Re[916]=-32'd9092; X_Re[84]=-32'd5662; X_Re[596]=32'd6326; X_Re[340]=-32'd4492; X_Re[852]=-32'd4310; X_Re[212]=-32'd6699; X_Re[724]=32'd3645; X_Re[468]=-32'd5322; X_Re[980]=32'd72; X_Re[52]=-32'd8022; X_Re[564]=-32'd10941; X_Re[308]=32'd21188; X_Re[820]=-32'd36128; X_Re[180]=32'd6839; X_Re[692]=32'd7248; X_Re[436]=-32'd1081; X_Re[948]=-32'd10342; X_Re[116]=-32'd5390; X_Re[628]=-32'd1703; X_Re[372]=-32'd9567; X_Re[884]=-32'd2829; X_Re[244]=-32'd1650; X_Re[756]=32'd33592; X_Re[500]=-32'd5174; X_Re[1012]=-32'd4157; X_Re[12]=-32'd4998; X_Re[524]=-32'd13655; X_Re[268]=-32'd12119; X_Re[780]=-32'd25781; X_Re[140]=-32'd36556; X_Re[652]=-32'd22939; X_Re[396]=32'd11030; X_Re[908]=32'd73677; X_Re[76]=32'd79471; X_Re[588]=-32'd12893; X_Re[332]=32'd45500; X_Re[844]=32'd22040; X_Re[204]=32'd113; X_Re[716]=32'd14818; X_Re[460]=32'd13157; X_Re[972]=32'd8849; X_Re[44]=32'd7302; X_Re[556]=32'd3742; X_Re[300]=32'd1597; X_Re[812]=-32'd4435; X_Re[172]=32'd12250; X_Re[684]=32'd14568; X_Re[428]=32'd5259; X_Re[940]=32'd6701; X_Re[108]=32'd1389; X_Re[620]=32'd5842; X_Re[364]=32'd4029; X_Re[876]=-32'd4858; X_Re[236]=-32'd3645; X_Re[748]=-32'd672; X_Re[492]=32'd4974; X_Re[1004]=32'd18305; X_Re[28]=32'd1586; X_Re[540]=32'd3644; X_Re[284]=-32'd3440; X_Re[796]=-32'd1443; X_Re[156]=32'd2725; X_Re[668]=-32'd1024; X_Re[412]=32'd5750; X_Re[924]=32'd2656; X_Re[92]=-32'd1000; X_Re[604]=-32'd3814; X_Re[348]=32'd12974; X_Re[860]=32'd444; X_Re[220]=-32'd135; X_Re[732]=-32'd17114; X_Re[476]=-32'd20408; X_Re[988]=32'd15575; X_Re[60]=32'd23887; X_Re[572]=-32'd5678; X_Re[316]=32'd2716; X_Re[828]=32'd7430; X_Re[188]=32'd5149; X_Re[700]=32'd1347; X_Re[444]=32'd198; X_Re[956]=32'd4325; X_Re[124]=32'd1647; X_Re[636]=32'd2362; X_Re[380]=-32'd4211; X_Re[892]=-32'd4557; X_Re[252]=32'd247; X_Re[764]=32'd561; X_Re[508]=-32'd2300; X_Re[1020]=-32'd2812; X_Re[2]=32'd4199; X_Re[514]=32'd6102; X_Re[258]=32'd2286; X_Re[770]=-32'd1321; X_Re[130]=32'd3711; X_Re[642]=-32'd4232; X_Re[386]=-32'd1814; X_Re[898]=-32'd1966; X_Re[66]=-32'd20260; X_Re[578]=-32'd12043; X_Re[322]=-32'd27418; X_Re[834]=32'd74501; X_Re[194]=-32'd12580; X_Re[706]=32'd51561; X_Re[450]=32'd38212; X_Re[962]=32'd5018; X_Re[34]=32'd10433; X_Re[546]=32'd1041; X_Re[290]=32'd4839; X_Re[802]=-32'd2275; X_Re[162]=32'd1240; X_Re[674]=-32'd9718; X_Re[418]=32'd19251; X_Re[930]=32'd15875; X_Re[98]=32'd24907; X_Re[610]=-32'd17830; X_Re[354]=32'd22972; X_Re[866]=-32'd15060; X_Re[226]=-32'd17454; X_Re[738]=32'd14979; X_Re[482]=32'd5478; X_Re[994]=32'd8163; X_Re[18]=32'd9653; X_Re[530]=32'd7815; X_Re[274]=-32'd4390; X_Re[786]=-32'd1107; X_Re[146]=32'd4921; X_Re[658]=32'd5641; X_Re[402]=32'd8048; X_Re[914]=32'd20142; X_Re[82]=32'd304; X_Re[594]=-32'd21717; X_Re[338]=-32'd15387; X_Re[850]=32'd910; X_Re[210]=-32'd5584; X_Re[722]=-32'd2360; X_Re[466]=-32'd4573; X_Re[978]=32'd4507; X_Re[50]=-32'd468; X_Re[562]=-32'd2353; X_Re[306]=-32'd4686; X_Re[818]=-32'd997; X_Re[178]=32'd3014; X_Re[690]=-32'd3343; X_Re[434]=-32'd10076; X_Re[946]=-32'd4711; X_Re[114]=-32'd119; X_Re[626]=-32'd8284; X_Re[370]=-32'd6385; X_Re[882]=32'd1001; X_Re[242]=-32'd20754; X_Re[754]=32'd6510; X_Re[498]=32'd9622; X_Re[1010]=-32'd12026; X_Re[10]=32'd2135; X_Re[522]=32'd4892; X_Re[266]=32'd14113; X_Re[778]=32'd12783; X_Re[138]=32'd9026; X_Re[650]=-32'd3351; X_Re[394]=-32'd3522; X_Re[906]=-32'd1883; X_Re[74]=-32'd2104; X_Re[586]=32'd2955; X_Re[330]=32'd1624; X_Re[842]=32'd9906; X_Re[202]=-32'd31088; X_Re[714]=-32'd69284; X_Re[458]=-32'd21741; X_Re[970]=32'd26174; X_Re[42]=32'd21107; X_Re[554]=32'd27095; X_Re[298]=32'd17744; X_Re[810]=32'd7843; X_Re[170]=32'd3575; X_Re[682]=32'd5268; X_Re[426]=32'd2275; X_Re[938]=32'd5093; X_Re[106]=32'd4152; X_Re[618]=32'd6587; X_Re[362]=32'd5706; X_Re[874]=32'd9694; X_Re[234]=-32'd219; X_Re[746]=-32'd6394; X_Re[490]=32'd9541; X_Re[1002]=32'd419; X_Re[26]=-32'd6571; X_Re[538]=-32'd12040; X_Re[282]=32'd12326; X_Re[794]=32'd13884; X_Re[154]=-32'd2894; X_Re[666]=32'd10079; X_Re[410]=32'd498; X_Re[922]=-32'd3106; X_Re[90]=32'd11603; X_Re[602]=-32'd2867; X_Re[346]=32'd3477; X_Re[858]=-32'd5876; X_Re[218]=-32'd3806; X_Re[730]=-32'd14665; X_Re[474]=32'd4292; X_Re[986]=32'd2298; X_Re[58]=32'd1134; X_Re[570]=32'd4562; X_Re[314]=-32'd4028; X_Re[826]=32'd1076; X_Re[186]=32'd1307; X_Re[698]=32'd1266; X_Re[442]=32'd5262; X_Re[954]=-32'd3120; X_Re[122]=32'd2932; X_Re[634]=32'd1223; X_Re[378]=32'd4195; X_Re[890]=32'd8723; X_Re[250]=32'd2828; X_Re[762]=-32'd2569; X_Re[506]=32'd185; X_Re[1018]=32'd791; X_Re[6]=32'd3287; X_Re[518]=32'd2779; X_Re[262]=32'd1264; X_Re[774]=32'd1993; X_Re[134]=-32'd2303; X_Re[646]=-32'd5224; X_Re[390]=32'd4668; X_Re[902]=-32'd484; X_Re[70]=-32'd1336; X_Re[582]=32'd3668; X_Re[326]=32'd7126; X_Re[838]=-32'd696; X_Re[198]=32'd5664; X_Re[710]=32'd6114; X_Re[454]=32'd5014; X_Re[966]=-32'd6974; X_Re[38]=32'd6777; X_Re[550]=-32'd5889; X_Re[294]=32'd8449; X_Re[806]=-32'd10760; X_Re[166]=-32'd14396; X_Re[678]=32'd3588; X_Re[422]=-32'd2938; X_Re[934]=32'd1930; X_Re[102]=32'd524; X_Re[614]=-32'd10544; X_Re[358]=-32'd1736; X_Re[870]=-32'd11328; X_Re[230]=32'd1017; X_Re[742]=-32'd2833; X_Re[486]=-32'd6321; X_Re[998]=-32'd7040; X_Re[22]=-32'd1046; X_Re[534]=-32'd4148; X_Re[278]=32'd8989; X_Re[790]=32'd14251; X_Re[150]=32'd1665; X_Re[662]=32'd9134; X_Re[406]=-32'd3527; X_Re[918]=32'd487; X_Re[86]=-32'd8390; X_Re[598]=-32'd7080; X_Re[342]=-32'd1364; X_Re[854]=-32'd5337; X_Re[214]=-32'd3161; X_Re[726]=32'd4474; X_Re[470]=32'd771; X_Re[982]=32'd11294; X_Re[54]=32'd710; X_Re[566]=32'd4136; X_Re[310]=-32'd1406; X_Re[822]=32'd1701; X_Re[182]=32'd3648; X_Re[694]=-32'd2515; X_Re[438]=32'd5600; X_Re[950]=-32'd1077; X_Re[118]=-32'd5290; X_Re[630]=-32'd1696; X_Re[374]=32'd253; X_Re[886]=-32'd3289; X_Re[246]=-32'd3339; X_Re[758]=32'd2039; X_Re[502]=-32'd239; X_Re[1014]=-32'd744; X_Re[14]=-32'd438; X_Re[526]=-32'd648; X_Re[270]=32'd4640; X_Re[782]=-32'd785; X_Re[142]=32'd3136; X_Re[654]=-32'd1347; X_Re[398]=-32'd2142; X_Re[910]=32'd81; X_Re[78]=-32'd610; X_Re[590]=32'd3765; X_Re[334]=32'd4386; X_Re[846]=32'd5782; X_Re[206]=-32'd4289; X_Re[718]=-32'd2578; X_Re[462]=-32'd7178; X_Re[974]=32'd2181; X_Re[46]=-32'd983; X_Re[558]=32'd478; X_Re[302]=-32'd12519; X_Re[814]=-32'd5800; X_Re[174]=-32'd11525; X_Re[686]=-32'd3360; X_Re[430]=-32'd9081; X_Re[942]=-32'd5005; X_Re[110]=32'd12347; X_Re[622]=32'd6589; X_Re[366]=-32'd4590; X_Re[878]=-32'd7421; X_Re[238]=-32'd7911; X_Re[750]=-32'd3481; X_Re[494]=32'd503; X_Re[1006]=-32'd4816; X_Re[30]=-32'd66; X_Re[542]=-32'd3201; X_Re[286]=-32'd4789; X_Re[798]=32'd468; X_Re[158]=32'd259; X_Re[670]=32'd2268; X_Re[414]=32'd14370; X_Re[926]=32'd7708; X_Re[94]=32'd12342; X_Re[606]=-32'd582; X_Re[350]=32'd3663; X_Re[862]=-32'd3903; X_Re[222]=-32'd8920; X_Re[734]=-32'd857; X_Re[478]=-32'd4053; X_Re[990]=-32'd1268; X_Re[62]=32'd5599; X_Re[574]=32'd3546; X_Re[318]=-32'd1949; X_Re[830]=-32'd2754; X_Re[190]=32'd5736; X_Re[702]=32'd725; X_Re[446]=-32'd6801; X_Re[958]=32'd4936; X_Re[126]=-32'd1656; X_Re[638]=-32'd1849; X_Re[382]=-32'd7295; X_Re[894]=32'd7049; X_Re[254]=-32'd804; X_Re[766]=32'd3487; X_Re[510]=-32'd2807; X_Re[1022]=32'd1575; X_Re[1]=-32'd1627; X_Re[513]=32'd1575; X_Re[257]=-32'd2807; X_Re[769]=32'd3487; X_Re[129]=-32'd804; X_Re[641]=32'd7049; X_Re[385]=-32'd7295; X_Re[897]=-32'd1849; X_Re[65]=-32'd1656; X_Re[577]=32'd4936; X_Re[321]=-32'd6801; X_Re[833]=32'd725; X_Re[193]=32'd5736; X_Re[705]=-32'd2754; X_Re[449]=-32'd1949; X_Re[961]=32'd3546; X_Re[33]=32'd5599; X_Re[545]=-32'd1268; X_Re[289]=-32'd4053; X_Re[801]=-32'd857; X_Re[161]=-32'd8920; X_Re[673]=-32'd3903; X_Re[417]=32'd3663; X_Re[929]=-32'd582; X_Re[97]=32'd12342; X_Re[609]=32'd7708; X_Re[353]=32'd14370; X_Re[865]=32'd2268; X_Re[225]=32'd259; X_Re[737]=32'd468; X_Re[481]=-32'd4789; X_Re[993]=-32'd3201; X_Re[17]=-32'd66; X_Re[529]=-32'd4816; X_Re[273]=32'd503; X_Re[785]=-32'd3481; X_Re[145]=-32'd7911; X_Re[657]=-32'd7421; X_Re[401]=-32'd4590; X_Re[913]=32'd6589; X_Re[81]=32'd12347; X_Re[593]=-32'd5005; X_Re[337]=-32'd9081; X_Re[849]=-32'd3360; X_Re[209]=-32'd11525; X_Re[721]=-32'd5800; X_Re[465]=-32'd12519; X_Re[977]=32'd478; X_Re[49]=-32'd983; X_Re[561]=32'd2181; X_Re[305]=-32'd7178; X_Re[817]=-32'd2578; X_Re[177]=-32'd4289; X_Re[689]=32'd5782; X_Re[433]=32'd4386; X_Re[945]=32'd3765; X_Re[113]=-32'd610; X_Re[625]=32'd81; X_Re[369]=-32'd2142; X_Re[881]=-32'd1347; X_Re[241]=32'd3136; X_Re[753]=-32'd785; X_Re[497]=32'd4640; X_Re[1009]=-32'd648; X_Re[9]=-32'd438; X_Re[521]=-32'd744; X_Re[265]=-32'd239; X_Re[777]=32'd2039; X_Re[137]=-32'd3339; X_Re[649]=-32'd3289; X_Re[393]=32'd253; X_Re[905]=-32'd1696; X_Re[73]=-32'd5290; X_Re[585]=-32'd1077; X_Re[329]=32'd5600; X_Re[841]=-32'd2515; X_Re[201]=32'd3648; X_Re[713]=32'd1701; X_Re[457]=-32'd1406; X_Re[969]=32'd4136; X_Re[41]=32'd710; X_Re[553]=32'd11294; X_Re[297]=32'd771; X_Re[809]=32'd4474; X_Re[169]=-32'd3161; X_Re[681]=-32'd5337; X_Re[425]=-32'd1364; X_Re[937]=-32'd7080; X_Re[105]=-32'd8390; X_Re[617]=32'd487; X_Re[361]=-32'd3527; X_Re[873]=32'd9134; X_Re[233]=32'd1665; X_Re[745]=32'd14251; X_Re[489]=32'd8989; X_Re[1001]=-32'd4148; X_Re[25]=-32'd1046; X_Re[537]=-32'd7040; X_Re[281]=-32'd6321; X_Re[793]=-32'd2833; X_Re[153]=32'd1017; X_Re[665]=-32'd11328; X_Re[409]=-32'd1736; X_Re[921]=-32'd10544; X_Re[89]=32'd524; X_Re[601]=32'd1930; X_Re[345]=-32'd2938; X_Re[857]=32'd3588; X_Re[217]=-32'd14396; X_Re[729]=-32'd10760; X_Re[473]=32'd8449; X_Re[985]=-32'd5889; X_Re[57]=32'd6777; X_Re[569]=-32'd6974; X_Re[313]=32'd5014; X_Re[825]=32'd6114; X_Re[185]=32'd5664; X_Re[697]=-32'd696; X_Re[441]=32'd7126; X_Re[953]=32'd3668; X_Re[121]=-32'd1336; X_Re[633]=-32'd484; X_Re[377]=32'd4668; X_Re[889]=-32'd5224; X_Re[249]=-32'd2303; X_Re[761]=32'd1993; X_Re[505]=32'd1264; X_Re[1017]=32'd2779; X_Re[5]=32'd3287; X_Re[517]=32'd791; X_Re[261]=32'd185; X_Re[773]=-32'd2569; X_Re[133]=32'd2828; X_Re[645]=32'd8723; X_Re[389]=32'd4195; X_Re[901]=32'd1223; X_Re[69]=32'd2932; X_Re[581]=-32'd3120; X_Re[325]=32'd5262; X_Re[837]=32'd1266; X_Re[197]=32'd1307; X_Re[709]=32'd1076; X_Re[453]=-32'd4028; X_Re[965]=32'd4562; X_Re[37]=32'd1134; X_Re[549]=32'd2298; X_Re[293]=32'd4292; X_Re[805]=-32'd14665; X_Re[165]=-32'd3806; X_Re[677]=-32'd5876; X_Re[421]=32'd3477; X_Re[933]=-32'd2867; X_Re[101]=32'd11603; X_Re[613]=-32'd3106; X_Re[357]=32'd498; X_Re[869]=32'd10079; X_Re[229]=-32'd2894; X_Re[741]=32'd13884; X_Re[485]=32'd12326; X_Re[997]=-32'd12040; X_Re[21]=-32'd6571; X_Re[533]=32'd419; X_Re[277]=32'd9541; X_Re[789]=-32'd6394; X_Re[149]=-32'd219; X_Re[661]=32'd9694; X_Re[405]=32'd5706; X_Re[917]=32'd6587; X_Re[85]=32'd4152; X_Re[597]=32'd5093; X_Re[341]=32'd2275; X_Re[853]=32'd5268; X_Re[213]=32'd3575; X_Re[725]=32'd7843; X_Re[469]=32'd17744; X_Re[981]=32'd27095; X_Re[53]=32'd21107; X_Re[565]=32'd26174; X_Re[309]=-32'd21741; X_Re[821]=-32'd69284; X_Re[181]=-32'd31088; X_Re[693]=32'd9906; X_Re[437]=32'd1624; X_Re[949]=32'd2955; X_Re[117]=-32'd2104; X_Re[629]=-32'd1883; X_Re[373]=-32'd3522; X_Re[885]=-32'd3351; X_Re[245]=32'd9026; X_Re[757]=32'd12783; X_Re[501]=32'd14113; X_Re[1013]=32'd4892; X_Re[13]=32'd2135; X_Re[525]=-32'd12026; X_Re[269]=32'd9622; X_Re[781]=32'd6510; X_Re[141]=-32'd20754; X_Re[653]=32'd1001; X_Re[397]=-32'd6385; X_Re[909]=-32'd8284; X_Re[77]=-32'd119; X_Re[589]=-32'd4711; X_Re[333]=-32'd10076; X_Re[845]=-32'd3343; X_Re[205]=32'd3014; X_Re[717]=-32'd997; X_Re[461]=-32'd4686; X_Re[973]=-32'd2353; X_Re[45]=-32'd468; X_Re[557]=32'd4507; X_Re[301]=-32'd4573; X_Re[813]=-32'd2360; X_Re[173]=-32'd5584; X_Re[685]=32'd910; X_Re[429]=-32'd15387; X_Re[941]=-32'd21717; X_Re[109]=32'd304; X_Re[621]=32'd20142; X_Re[365]=32'd8048; X_Re[877]=32'd5641; X_Re[237]=32'd4921; X_Re[749]=-32'd1107; X_Re[493]=-32'd4390; X_Re[1005]=32'd7815; X_Re[29]=32'd9653; X_Re[541]=32'd8163; X_Re[285]=32'd5478; X_Re[797]=32'd14979; X_Re[157]=-32'd17454; X_Re[669]=-32'd15060; X_Re[413]=32'd22972; X_Re[925]=-32'd17830; X_Re[93]=32'd24907; X_Re[605]=32'd15875; X_Re[349]=32'd19251; X_Re[861]=-32'd9718; X_Re[221]=32'd1240; X_Re[733]=-32'd2275; X_Re[477]=32'd4839; X_Re[989]=32'd1041; X_Re[61]=32'd10433; X_Re[573]=32'd5018; X_Re[317]=32'd38212; X_Re[829]=32'd51561; X_Re[189]=-32'd12580; X_Re[701]=32'd74501; X_Re[445]=-32'd27418; X_Re[957]=-32'd12043; X_Re[125]=-32'd20260; X_Re[637]=-32'd1966; X_Re[381]=-32'd1814; X_Re[893]=-32'd4232; X_Re[253]=32'd3711; X_Re[765]=-32'd1321; X_Re[509]=32'd2286; X_Re[1021]=32'd6102; X_Re[3]=32'd4199; X_Re[515]=-32'd2812; X_Re[259]=-32'd2300; X_Re[771]=32'd561; X_Re[131]=32'd247; X_Re[643]=-32'd4557; X_Re[387]=-32'd4211; X_Re[899]=32'd2362; X_Re[67]=32'd1647; X_Re[579]=32'd4325; X_Re[323]=32'd198; X_Re[835]=32'd1347; X_Re[195]=32'd5149; X_Re[707]=32'd7430; X_Re[451]=32'd2716; X_Re[963]=-32'd5678; X_Re[35]=32'd23887; X_Re[547]=32'd15575; X_Re[291]=-32'd20408; X_Re[803]=-32'd17114; X_Re[163]=-32'd135; X_Re[675]=32'd444; X_Re[419]=32'd12974; X_Re[931]=-32'd3814; X_Re[99]=-32'd1000; X_Re[611]=32'd2656; X_Re[355]=32'd5750; X_Re[867]=-32'd1024; X_Re[227]=32'd2725; X_Re[739]=-32'd1443; X_Re[483]=-32'd3440; X_Re[995]=32'd3644; X_Re[19]=32'd1586; X_Re[531]=32'd18305; X_Re[275]=32'd4974; X_Re[787]=-32'd672; X_Re[147]=-32'd3645; X_Re[659]=-32'd4858; X_Re[403]=32'd4029; X_Re[915]=32'd5842; X_Re[83]=32'd1389; X_Re[595]=32'd6701; X_Re[339]=32'd5259; X_Re[851]=32'd14568; X_Re[211]=32'd12250; X_Re[723]=-32'd4435; X_Re[467]=32'd1597; X_Re[979]=32'd3742; X_Re[51]=32'd7302; X_Re[563]=32'd8849; X_Re[307]=32'd13157; X_Re[819]=32'd14818; X_Re[179]=32'd113; X_Re[691]=32'd22040; X_Re[435]=32'd45500; X_Re[947]=-32'd12893; X_Re[115]=32'd79471; X_Re[627]=32'd73677; X_Re[371]=32'd11030; X_Re[883]=-32'd22939; X_Re[243]=-32'd36556; X_Re[755]=-32'd25781; X_Re[499]=-32'd12119; X_Re[1011]=-32'd13655; X_Re[11]=-32'd4998; X_Re[523]=-32'd4157; X_Re[267]=-32'd5174; X_Re[779]=32'd33592; X_Re[139]=-32'd1650; X_Re[651]=-32'd2829; X_Re[395]=-32'd9567; X_Re[907]=-32'd1703; X_Re[75]=-32'd5390; X_Re[587]=-32'd10342; X_Re[331]=-32'd1081; X_Re[843]=32'd7248; X_Re[203]=32'd6839; X_Re[715]=-32'd36128; X_Re[459]=32'd21188; X_Re[971]=-32'd10941; X_Re[43]=-32'd8022; X_Re[555]=32'd72; X_Re[299]=-32'd5322; X_Re[811]=32'd3645; X_Re[171]=-32'd6699; X_Re[683]=-32'd4310; X_Re[427]=-32'd4492; X_Re[939]=32'd6326; X_Re[107]=-32'd5662; X_Re[619]=-32'd9092; X_Re[363]=32'd2843; X_Re[875]=-32'd7142; X_Re[235]=-32'd18047; X_Re[747]=32'd7595; X_Re[491]=-32'd13945; X_Re[1003]=-32'd53731; X_Re[27]=32'd44207; X_Re[539]=-32'd26098; X_Re[283]=32'd43192; X_Re[795]=32'd16551; X_Re[155]=-32'd9583; X_Re[667]=32'd7908; X_Re[411]=-32'd785; X_Re[923]=32'd5927; X_Re[91]=32'd4481; X_Re[603]=32'd9251; X_Re[347]=32'd8099; X_Re[859]=32'd3541; X_Re[219]=32'd1191; X_Re[731]=32'd5648; X_Re[475]=32'd7001; X_Re[987]=32'd1621; X_Re[59]=32'd2346; X_Re[571]=-32'd7572; X_Re[315]=32'd8862; X_Re[827]=32'd24684; X_Re[187]=-32'd14770; X_Re[699]=-32'd7719; X_Re[443]=-32'd2938; X_Re[955]=-32'd10221; X_Re[123]=32'd4423; X_Re[635]=-32'd59599; X_Re[379]=32'd70108; X_Re[891]=32'd348596; X_Re[251]=32'd28921; X_Re[763]=-32'd5217; X_Re[507]=32'd1626; X_Re[1019]=-32'd5956; X_Re[7]=-32'd2026; X_Re[519]=-32'd2025; X_Re[263]=32'd242; X_Re[775]=32'd11710; X_Re[135]=-32'd653; X_Re[647]=32'd4346; X_Re[391]=32'd16199; X_Re[903]=-32'd8956; X_Re[71]=32'd35868; X_Re[583]=-32'd93185; X_Re[327]=-32'd14034; X_Re[839]=32'd24008; X_Re[199]=32'd7848; X_Re[711]=32'd3472; X_Re[455]=32'd8206; X_Re[967]=32'd4331; X_Re[39]=-32'd4449; X_Re[551]=32'd7264; X_Re[295]=-32'd870; X_Re[807]=32'd13462; X_Re[167]=32'd2968; X_Re[679]=32'd20766; X_Re[423]=32'd36890; X_Re[935]=-32'd33732; X_Re[103]=-32'd8783; X_Re[615]=-32'd6999; X_Re[359]=-32'd429; X_Re[871]=32'd2850; X_Re[231]=32'd2743; X_Re[743]=32'd3784; X_Re[487]=-32'd6194; X_Re[999]=-32'd15483; X_Re[23]=-32'd1423; X_Re[535]=-32'd32083; X_Re[279]=32'd53368; X_Re[791]=32'd11635; X_Re[151]=32'd10361; X_Re[663]=32'd19519; X_Re[407]=32'd13322; X_Re[919]=32'd328; X_Re[87]=32'd12647; X_Re[599]=32'd6553; X_Re[343]=32'd508; X_Re[855]=32'd1599; X_Re[215]=32'd7487; X_Re[727]=32'd10478; X_Re[471]=32'd5014; X_Re[983]=32'd21865; X_Re[55]=-32'd103143; X_Re[567]=-32'd322659; X_Re[311]=-32'd2159; X_Re[823]=32'd18835; X_Re[183]=32'd15514; X_Re[695]=32'd20953; X_Re[439]=32'd24094; X_Re[951]=32'd27560; X_Re[119]=32'd20529; X_Re[631]=32'd86424; X_Re[375]=32'd24689; X_Re[887]=32'd98286; X_Re[247]=32'd25897; X_Re[759]=-32'd220475; X_Re[503]=-32'd350559; X_Re[1015]=-32'd84078; X_Re[15]=-32'd89550; X_Re[527]=-32'd73725; X_Re[271]=-32'd68355; X_Re[783]=-32'd76563; X_Re[143]=-32'd374488; X_Re[655]=32'd172680; X_Re[399]=32'd99801; X_Re[911]=32'd16164; X_Re[79]=32'd19028; X_Re[591]=-32'd2465; X_Re[335]=-32'd32042; X_Re[847]=32'd200812; X_Re[207]=32'd3041; X_Re[719]=32'd44296; X_Re[463]=32'd18707; X_Re[975]=32'd19509; X_Re[47]=32'd37484; X_Re[559]=32'd35091; X_Re[303]=32'd7926; X_Re[815]=32'd32371; X_Re[175]=32'd71278; X_Re[687]=32'd19080; X_Re[431]=32'd48085; X_Re[943]=32'd77266; X_Re[111]=32'd422815; X_Re[623]=-32'd219111; X_Re[367]=-32'd92155; X_Re[879]=-32'd33674; X_Re[239]=-32'd57943; X_Re[751]=32'd31774; X_Re[495]=-32'd22086; X_Re[1007]=-32'd10798; X_Re[31]=-32'd20014; X_Re[543]=-32'd23713; X_Re[287]=-32'd38433; X_Re[799]=-32'd23890; X_Re[159]=-32'd34797; X_Re[671]=-32'd73347; X_Re[415]=32'd41646; X_Re[927]=32'd2592; X_Re[95]=-32'd5577; X_Re[607]=32'd13800; X_Re[351]=-32'd4748; X_Re[863]=-32'd19342; X_Re[223]=32'd1037; X_Re[735]=-32'd54871; X_Re[479]=-32'd32079; X_Re[991]=32'd41019; X_Re[63]=-32'd12426; X_Re[575]=32'd16013; X_Re[319]=32'd2080; X_Re[831]=-32'd40016; X_Re[191]=-32'd7187; X_Re[703]=32'd71943; X_Re[447]=-32'd45666; X_Re[959]=-32'd166613; X_Re[127]=-32'd5662; X_Re[639]=-32'd45742; X_Re[383]=-32'd13493; X_Re[895]=-32'd8097; X_Re[255]=-32'd3178; X_Re[767]=-32'd3237; X_Re[511]=32'd8055; X_Re[1023]=32'd3344; 
		X_Im[0]=32'd0; X_Im[512]=-32'd1486; X_Im[256]=-32'd12913; X_Im[768]=-32'd28663; X_Im[128]=-32'd30790; X_Im[640]=-32'd34136; X_Im[384]=-32'd73376; X_Im[896]=32'd48603; X_Im[64]=-32'd40194; X_Im[576]=32'd139265; X_Im[320]=32'd35545; X_Im[832]=32'd12968; X_Im[192]=32'd25657; X_Im[704]=32'd94271; X_Im[448]=-32'd12300; X_Im[960]=32'd15022; X_Im[32]=32'd6583; X_Im[544]=32'd4976; X_Im[288]=32'd64934; X_Im[800]=32'd42162; X_Im[160]=32'd46940; X_Im[672]=32'd19111; X_Im[416]=32'd21141; X_Im[928]=-32'd17590; X_Im[96]=32'd12985; X_Im[608]=32'd8041; X_Im[352]=-32'd11679; X_Im[864]=32'd20701; X_Im[224]=32'd28244; X_Im[736]=32'd25853; X_Im[480]=32'd31296; X_Im[992]=32'd36200; X_Im[16]=32'd37022; X_Im[528]=32'd46075; X_Im[272]=32'd52457; X_Im[784]=32'd88522; X_Im[144]=32'd67934; X_Im[656]=32'd87548; X_Im[400]=32'd154365; X_Im[912]=32'd611736; X_Im[80]=-32'd332002; X_Im[592]=-32'd114939; X_Im[336]=-32'd77472; X_Im[848]=-32'd66258; X_Im[208]=-32'd22530; X_Im[720]=32'd40748; X_Im[464]=-32'd5987; X_Im[976]=32'd85512; X_Im[48]=-32'd26484; X_Im[560]=-32'd30607; X_Im[304]=-32'd7730; X_Im[816]=-32'd22785; X_Im[176]=32'd11192; X_Im[688]=32'd87188; X_Im[432]=-32'd32459; X_Im[944]=-32'd34272; X_Im[112]=-32'd44533; X_Im[624]=-32'd4368; X_Im[368]=-32'd88372; X_Im[880]=-32'd182053; X_Im[240]=32'd6643; X_Im[752]=-32'd5077; X_Im[496]=32'd8026; X_Im[1008]=32'd4488; X_Im[8]=-32'd10776; X_Im[520]=32'd6967; X_Im[264]=32'd124522; X_Im[776]=-32'd714901; X_Im[136]=32'd151433; X_Im[648]=32'd4696; X_Im[392]=32'd1668; X_Im[904]=-32'd63305; X_Im[72]=-32'd55297; X_Im[584]=-32'd10093; X_Im[328]=-32'd22629; X_Im[840]=-32'd33190; X_Im[200]=-32'd27931; X_Im[712]=-32'd40605; X_Im[456]=-32'd64712; X_Im[968]=-32'd183414; X_Im[40]=32'd70691; X_Im[552]=32'd75688; X_Im[296]=32'd34833; X_Im[808]=32'd23195; X_Im[168]=32'd12639; X_Im[680]=32'd14039; X_Im[424]=32'd9496; X_Im[936]=32'd11844; X_Im[104]=32'd46374; X_Im[616]=32'd66525; X_Im[360]=-32'd34823; X_Im[872]=-32'd30190; X_Im[232]=-32'd24689; X_Im[744]=-32'd7105; X_Im[488]=-32'd25124; X_Im[1000]=-32'd1563; X_Im[24]=-32'd11538; X_Im[536]=-32'd1057; X_Im[280]=32'd6873; X_Im[792]=-32'd1126; X_Im[152]=32'd2601; X_Im[664]=-32'd991; X_Im[408]=-32'd8961; X_Im[920]=-32'd5380; X_Im[88]=-32'd21730; X_Im[600]=-32'd11776; X_Im[344]=32'd22830; X_Im[856]=32'd8519; X_Im[216]=32'd4870; X_Im[728]=-32'd5188; X_Im[472]=-32'd8343; X_Im[984]=-32'd2572; X_Im[56]=-32'd32539; X_Im[568]=-32'd15082; X_Im[312]=-32'd32568; X_Im[824]=-32'd32225; X_Im[184]=-32'd54085; X_Im[696]=-32'd114821; X_Im[440]=-32'd30338; X_Im[952]=32'd133139; X_Im[120]=32'd159144; X_Im[632]=32'd4768; X_Im[376]=32'd32457; X_Im[888]=32'd8339; X_Im[248]=32'd21897; X_Im[760]=32'd22138; X_Im[504]=32'd17927; X_Im[1016]=32'd16925; X_Im[4]=32'd14000; X_Im[516]=32'd18947; X_Im[260]=32'd24502; X_Im[772]=32'd43848; X_Im[132]=32'd77885; X_Im[644]=-32'd29326; X_Im[388]=-32'd175459; X_Im[900]=32'd148481; X_Im[68]=-32'd17815; X_Im[580]=32'd13203; X_Im[324]=32'd5862; X_Im[836]=32'd9077; X_Im[196]=32'd17405; X_Im[708]=32'd42849; X_Im[452]=32'd10751; X_Im[964]=32'd7477; X_Im[36]=-32'd5964; X_Im[548]=32'd1260; X_Im[292]=32'd1; X_Im[804]=-32'd1974; X_Im[164]=-32'd339; X_Im[676]=32'd766; X_Im[420]=32'd3011; X_Im[932]=32'd4257; X_Im[100]=-32'd2636; X_Im[612]=32'd5153; X_Im[356]=-32'd89; X_Im[868]=-32'd676; X_Im[228]=-32'd4537; X_Im[740]=-32'd25667; X_Im[484]=-32'd38556; X_Im[996]=32'd73732; X_Im[20]=-32'd30401; X_Im[532]=-32'd45472; X_Im[276]=32'd10007; X_Im[788]=32'd3204; X_Im[148]=32'd14901; X_Im[660]=32'd8129; X_Im[404]=32'd9738; X_Im[916]=32'd5613; X_Im[84]=32'd7049; X_Im[596]=-32'd3376; X_Im[340]=32'd8437; X_Im[852]=-32'd3625; X_Im[212]=32'd5402; X_Im[724]=32'd6524; X_Im[468]=-32'd1992; X_Im[980]=32'd686; X_Im[52]=32'd2011; X_Im[564]=32'd10031; X_Im[308]=-32'd17162; X_Im[820]=32'd19053; X_Im[180]=32'd13251; X_Im[692]=32'd1537; X_Im[436]=-32'd2780; X_Im[948]=32'd1474; X_Im[116]=32'd11040; X_Im[628]=-32'd1846; X_Im[372]=32'd2570; X_Im[884]=32'd25003; X_Im[244]=32'd11756; X_Im[756]=-32'd15558; X_Im[500]=32'd4871; X_Im[1012]=32'd10858; X_Im[12]=32'd1345; X_Im[524]=32'd16888; X_Im[268]=32'd12192; X_Im[780]=32'd22139; X_Im[140]=32'd30560; X_Im[652]=32'd64467; X_Im[396]=32'd98891; X_Im[908]=32'd63798; X_Im[76]=32'd58461; X_Im[588]=-32'd134452; X_Im[332]=32'd4902; X_Im[844]=-32'd37908; X_Im[204]=-32'd25585; X_Im[716]=-32'd13828; X_Im[460]=-32'd20123; X_Im[972]=-32'd19440; X_Im[44]=-32'd13366; X_Im[556]=-32'd11450; X_Im[300]=-32'd10890; X_Im[812]=-32'd11523; X_Im[172]=32'd1116; X_Im[684]=-32'd18114; X_Im[428]=-32'd11902; X_Im[940]=-32'd12952; X_Im[108]=-32'd7149; X_Im[620]=-32'd13536; X_Im[364]=-32'd12617; X_Im[876]=-32'd10742; X_Im[236]=-32'd5421; X_Im[748]=-32'd6244; X_Im[492]=32'd9592; X_Im[1004]=-32'd11491; X_Im[28]=-32'd1015; X_Im[540]=-32'd7961; X_Im[284]=-32'd7358; X_Im[796]=-32'd4288; X_Im[156]=-32'd1380; X_Im[668]=32'd759; X_Im[412]=-32'd647; X_Im[924]=-32'd1958; X_Im[92]=-32'd4480; X_Im[604]=-32'd11132; X_Im[348]=-32'd3671; X_Im[860]=-32'd15006; X_Im[220]=32'd2644; X_Im[732]=-32'd16467; X_Im[476]=-32'd5439; X_Im[988]=-32'd7724; X_Im[60]=-32'd5725; X_Im[572]=-32'd3686; X_Im[316]=32'd15040; X_Im[828]=32'd543; X_Im[188]=-32'd2579; X_Im[700]=-32'd4814; X_Im[444]=-32'd6068; X_Im[956]=32'd93; X_Im[124]=-32'd1652; X_Im[636]=-32'd4159; X_Im[380]=-32'd2390; X_Im[892]=-32'd2923; X_Im[252]=32'd3903; X_Im[764]=-32'd3797; X_Im[508]=32'd5393; X_Im[1020]=32'd7721; X_Im[2]=-32'd2824; X_Im[514]=32'd658; X_Im[258]=32'd4283; X_Im[770]=-32'd7941; X_Im[130]=32'd1441; X_Im[642]=-32'd1942; X_Im[386]=-32'd7979; X_Im[898]=-32'd12687; X_Im[66]=-32'd5325; X_Im[578]=32'd16399; X_Im[322]=32'd8936; X_Im[834]=32'd19877; X_Im[194]=-32'd21451; X_Im[706]=32'd67060; X_Im[450]=-32'd39729; X_Im[962]=-32'd13946; X_Im[34]=-32'd11436; X_Im[546]=-32'd10534; X_Im[290]=32'd5730; X_Im[802]=32'd2246; X_Im[162]=-32'd857; X_Im[674]=32'd10964; X_Im[418]=32'd4875; X_Im[930]=-32'd1199; X_Im[98]=-32'd14740; X_Im[610]=-32'd23781; X_Im[354]=32'd22921; X_Im[866]=-32'd29632; X_Im[226]=32'd2578; X_Im[738]=-32'd15490; X_Im[482]=-32'd5407; X_Im[994]=-32'd4612; X_Im[18]=-32'd9143; X_Im[530]=-32'd9133; X_Im[274]=-32'd13702; X_Im[786]=-32'd2488; X_Im[146]=-32'd10580; X_Im[658]=32'd3262; X_Im[402]=-32'd6800; X_Im[914]=-32'd11007; X_Im[82]=-32'd39175; X_Im[594]=32'd1411; X_Im[338]=32'd21317; X_Im[850]=32'd2085; X_Im[210]=32'd412; X_Im[722]=-32'd3416; X_Im[466]=32'd3541; X_Im[978]=-32'd7040; X_Im[50]=-32'd2408; X_Im[562]=-32'd4202; X_Im[306]=-32'd6966; X_Im[818]=-32'd7091; X_Im[178]=-32'd4959; X_Im[690]=-32'd12769; X_Im[434]=-32'd2306; X_Im[946]=-32'd1316; X_Im[114]=32'd372; X_Im[626]=32'd1369; X_Im[370]=32'd4235; X_Im[882]=32'd5924; X_Im[242]=32'd1375; X_Im[754]=32'd2672; X_Im[498]=32'd17029; X_Im[1010]=-32'd8068; X_Im[10]=-32'd6176; X_Im[522]=-32'd5513; X_Im[266]=-32'd15716; X_Im[778]=32'd17029; X_Im[138]=32'd7765; X_Im[650]=-32'd1706; X_Im[394]=32'd3634; X_Im[906]=-32'd2045; X_Im[74]=-32'd3852; X_Im[586]=-32'd3748; X_Im[330]=32'd7865; X_Im[842]=32'd1947; X_Im[202]=32'd5505; X_Im[714]=32'd5105; X_Im[458]=32'd51981; X_Im[970]=32'd13172; X_Im[42]=-32'd8142; X_Im[554]=-32'd16513; X_Im[298]=-32'd5668; X_Im[810]=-32'd10835; X_Im[170]=-32'd7954; X_Im[682]=32'd983; X_Im[426]=-32'd2868; X_Im[938]=-32'd3944; X_Im[106]=-32'd2702; X_Im[618]=-32'd4609; X_Im[362]=-32'd1238; X_Im[874]=32'd1182; X_Im[234]=-32'd4593; X_Im[746]=-32'd648; X_Im[490]=-32'd2063; X_Im[1002]=-32'd7577; X_Im[26]=32'd740; X_Im[538]=-32'd5182; X_Im[282]=32'd2008; X_Im[794]=32'd2692; X_Im[154]=32'd8843; X_Im[666]=32'd13482; X_Im[410]=-32'd6697; X_Im[922]=32'd532; X_Im[90]=32'd13; X_Im[602]=32'd3253; X_Im[346]=-32'd6839; X_Im[858]=32'd2645; X_Im[218]=-32'd14516; X_Im[730]=-32'd3828; X_Im[474]=-32'd5213; X_Im[986]=-32'd1412; X_Im[58]=-32'd5540; X_Im[570]=-32'd3715; X_Im[314]=-32'd7968; X_Im[826]=-32'd3156; X_Im[186]=-32'd6089; X_Im[698]=32'd305; X_Im[442]=32'd1943; X_Im[954]=-32'd22; X_Im[122]=-32'd2067; X_Im[634]=-32'd4206; X_Im[378]=-32'd8335; X_Im[890]=-32'd4071; X_Im[250]=-32'd3027; X_Im[762]=-32'd4207; X_Im[506]=32'd3024; X_Im[1018]=-32'd1894; X_Im[6]=-32'd198; X_Im[518]=-32'd1914; X_Im[262]=-32'd3905; X_Im[774]=-32'd1740; X_Im[134]=-32'd4085; X_Im[646]=-32'd4159; X_Im[390]=32'd6551; X_Im[902]=-32'd1969; X_Im[70]=32'd629; X_Im[582]=-32'd183; X_Im[326]=32'd2484; X_Im[838]=32'd4080; X_Im[198]=-32'd6235; X_Im[710]=32'd4880; X_Im[454]=32'd757; X_Im[966]=-32'd4999; X_Im[38]=32'd654; X_Im[550]=-32'd15284; X_Im[294]=-32'd12873; X_Im[806]=-32'd18119; X_Im[166]=32'd2731; X_Im[678]=-32'd5999; X_Im[422]=-32'd5323; X_Im[934]=-32'd4532; X_Im[102]=-32'd10189; X_Im[614]=-32'd6429; X_Im[358]=-32'd1661; X_Im[870]=-32'd5113; X_Im[230]=32'd4613; X_Im[742]=-32'd1782; X_Im[486]=-32'd4460; X_Im[998]=32'd1253; X_Im[22]=32'd2230; X_Im[534]=32'd6426; X_Im[278]=32'd1246; X_Im[790]=-32'd3504; X_Im[150]=-32'd9277; X_Im[662]=-32'd4114; X_Im[406]=-32'd1129; X_Im[918]=-32'd5825; X_Im[86]=-32'd563; X_Im[598]=32'd6218; X_Im[342]=-32'd1591; X_Im[854]=32'd6354; X_Im[214]=32'd7503; X_Im[726]=-32'd7132; X_Im[470]=-32'd8735; X_Im[982]=-32'd5977; X_Im[54]=32'd5753; X_Im[566]=-32'd5444; X_Im[310]=-32'd802; X_Im[822]=-32'd1534; X_Im[182]=32'd8611; X_Im[694]=-32'd983; X_Im[438]=32'd1747; X_Im[950]=-32'd2351; X_Im[118]=-32'd5723; X_Im[630]=-32'd411; X_Im[374]=-32'd5597; X_Im[886]=32'd5090; X_Im[246]=32'd6770; X_Im[758]=-32'd555; X_Im[502]=-32'd3432; X_Im[1014]=-32'd277; X_Im[14]=-32'd2007; X_Im[526]=-32'd922; X_Im[270]=32'd1828; X_Im[782]=-32'd623; X_Im[142]=-32'd3972; X_Im[654]=-32'd4785; X_Im[398]=-32'd376; X_Im[910]=32'd1659; X_Im[78]=-32'd261; X_Im[590]=-32'd1479; X_Im[334]=-32'd2322; X_Im[846]=-32'd5757; X_Im[206]=-32'd10124; X_Im[718]=-32'd979; X_Im[462]=32'd8593; X_Im[974]=-32'd4476; X_Im[46]=-32'd7906; X_Im[558]=-32'd15385; X_Im[302]=-32'd12030; X_Im[814]=-32'd4084; X_Im[174]=-32'd605; X_Im[686]=32'd5764; X_Im[430]=-32'd17361; X_Im[942]=-32'd64; X_Im[110]=32'd3406; X_Im[622]=32'd2153; X_Im[366]=-32'd3854; X_Im[878]=32'd5348; X_Im[238]=32'd9053; X_Im[750]=-32'd5211; X_Im[494]=32'd4238; X_Im[1006]=32'd2016; X_Im[30]=-32'd1592; X_Im[542]=32'd3580; X_Im[286]=32'd7527; X_Im[798]=32'd1098; X_Im[158]=32'd4156; X_Im[670]=32'd2445; X_Im[414]=-32'd8454; X_Im[926]=-32'd493; X_Im[94]=32'd2760; X_Im[606]=-32'd12007; X_Im[350]=-32'd1216; X_Im[862]=-32'd982; X_Im[222]=-32'd7836; X_Im[734]=32'd6778; X_Im[478]=-32'd2138; X_Im[990]=32'd2606; X_Im[62]=-32'd7651; X_Im[574]=32'd15514; X_Im[318]=-32'd1274; X_Im[830]=32'd7193; X_Im[190]=-32'd3310; X_Im[702]=-32'd2899; X_Im[446]=32'd5410; X_Im[958]=32'd2766; X_Im[126]=-32'd5843; X_Im[638]=-32'd5049; X_Im[382]=-32'd192; X_Im[894]=32'd4135; X_Im[254]=-32'd5963; X_Im[766]=-32'd4336; X_Im[510]=32'd2465; X_Im[1022]=-32'd1617; X_Im[1]=32'd0; X_Im[513]=32'd1617; X_Im[257]=-32'd2465; X_Im[769]=32'd4336; X_Im[129]=32'd5963; X_Im[641]=-32'd4135; X_Im[385]=32'd192; X_Im[897]=32'd5049; X_Im[65]=32'd5843; X_Im[577]=-32'd2766; X_Im[321]=-32'd5410; X_Im[833]=32'd2899; X_Im[193]=32'd3310; X_Im[705]=-32'd7193; X_Im[449]=32'd1274; X_Im[961]=-32'd15514; X_Im[33]=32'd7651; X_Im[545]=-32'd2606; X_Im[289]=32'd2138; X_Im[801]=-32'd6778; X_Im[161]=32'd7836; X_Im[673]=32'd982; X_Im[417]=32'd1216; X_Im[929]=32'd12007; X_Im[97]=-32'd2760; X_Im[609]=32'd493; X_Im[353]=32'd8454; X_Im[865]=-32'd2445; X_Im[225]=-32'd4156; X_Im[737]=-32'd1098; X_Im[481]=-32'd7527; X_Im[993]=-32'd3580; X_Im[17]=32'd1592; X_Im[529]=-32'd2016; X_Im[273]=-32'd4238; X_Im[785]=32'd5211; X_Im[145]=-32'd9053; X_Im[657]=-32'd5348; X_Im[401]=32'd3854; X_Im[913]=-32'd2153; X_Im[81]=-32'd3406; X_Im[593]=32'd64; X_Im[337]=32'd17361; X_Im[849]=-32'd5764; X_Im[209]=32'd605; X_Im[721]=32'd4084; X_Im[465]=32'd12030; X_Im[977]=32'd15385; X_Im[49]=32'd7906; X_Im[561]=32'd4476; X_Im[305]=-32'd8593; X_Im[817]=32'd979; X_Im[177]=32'd10124; X_Im[689]=32'd5757; X_Im[433]=32'd2322; X_Im[945]=32'd1479; X_Im[113]=32'd261; X_Im[625]=-32'd1659; X_Im[369]=32'd376; X_Im[881]=32'd4785; X_Im[241]=32'd3972; X_Im[753]=32'd623; X_Im[497]=-32'd1828; X_Im[1009]=32'd922; X_Im[9]=32'd2007; X_Im[521]=32'd277; X_Im[265]=32'd3432; X_Im[777]=32'd555; X_Im[137]=-32'd6770; X_Im[649]=-32'd5090; X_Im[393]=32'd5597; X_Im[905]=32'd411; X_Im[73]=32'd5723; X_Im[585]=32'd2351; X_Im[329]=-32'd1747; X_Im[841]=32'd983; X_Im[201]=-32'd8611; X_Im[713]=32'd1534; X_Im[457]=32'd802; X_Im[969]=32'd5444; X_Im[41]=-32'd5753; X_Im[553]=32'd5977; X_Im[297]=32'd8735; X_Im[809]=32'd7132; X_Im[169]=-32'd7503; X_Im[681]=-32'd6354; X_Im[425]=32'd1591; X_Im[937]=-32'd6218; X_Im[105]=32'd563; X_Im[617]=32'd5825; X_Im[361]=32'd1129; X_Im[873]=32'd4114; X_Im[233]=32'd9277; X_Im[745]=32'd3504; X_Im[489]=-32'd1246; X_Im[1001]=-32'd6426; X_Im[25]=-32'd2230; X_Im[537]=-32'd1253; X_Im[281]=32'd4460; X_Im[793]=32'd1782; X_Im[153]=-32'd4613; X_Im[665]=32'd5113; X_Im[409]=32'd1661; X_Im[921]=32'd6429; X_Im[89]=32'd10189; X_Im[601]=32'd4532; X_Im[345]=32'd5323; X_Im[857]=32'd5999; X_Im[217]=-32'd2731; X_Im[729]=32'd18119; X_Im[473]=32'd12873; X_Im[985]=32'd15284; X_Im[57]=-32'd654; X_Im[569]=32'd4999; X_Im[313]=-32'd757; X_Im[825]=-32'd4880; X_Im[185]=32'd6235; X_Im[697]=-32'd4080; X_Im[441]=-32'd2484; X_Im[953]=32'd183; X_Im[121]=-32'd629; X_Im[633]=32'd1969; X_Im[377]=-32'd6551; X_Im[889]=32'd4159; X_Im[249]=32'd4085; X_Im[761]=32'd1740; X_Im[505]=32'd3905; X_Im[1017]=32'd1914; X_Im[5]=32'd198; X_Im[517]=32'd1894; X_Im[261]=-32'd3024; X_Im[773]=32'd4207; X_Im[133]=32'd3027; X_Im[645]=32'd4071; X_Im[389]=32'd8335; X_Im[901]=32'd4206; X_Im[69]=32'd2067; X_Im[581]=32'd22; X_Im[325]=-32'd1943; X_Im[837]=-32'd305; X_Im[197]=32'd6089; X_Im[709]=32'd3156; X_Im[453]=32'd7968; X_Im[965]=32'd3715; X_Im[37]=32'd5540; X_Im[549]=32'd1412; X_Im[293]=32'd5213; X_Im[805]=32'd3828; X_Im[165]=32'd14516; X_Im[677]=-32'd2645; X_Im[421]=32'd6839; X_Im[933]=-32'd3253; X_Im[101]=-32'd13; X_Im[613]=-32'd532; X_Im[357]=32'd6697; X_Im[869]=-32'd13482; X_Im[229]=-32'd8843; X_Im[741]=-32'd2692; X_Im[485]=-32'd2008; X_Im[997]=32'd5182; X_Im[21]=-32'd740; X_Im[533]=32'd7577; X_Im[277]=32'd2063; X_Im[789]=32'd648; X_Im[149]=32'd4593; X_Im[661]=-32'd1182; X_Im[405]=32'd1238; X_Im[917]=32'd4609; X_Im[85]=32'd2702; X_Im[597]=32'd3944; X_Im[341]=32'd2868; X_Im[853]=-32'd983; X_Im[213]=32'd7954; X_Im[725]=32'd10835; X_Im[469]=32'd5668; X_Im[981]=32'd16513; X_Im[53]=32'd8142; X_Im[565]=-32'd13172; X_Im[309]=-32'd51981; X_Im[821]=-32'd5105; X_Im[181]=-32'd5505; X_Im[693]=-32'd1947; X_Im[437]=-32'd7865; X_Im[949]=32'd3748; X_Im[117]=32'd3852; X_Im[629]=32'd2045; X_Im[373]=-32'd3634; X_Im[885]=32'd1706; X_Im[245]=-32'd7765; X_Im[757]=-32'd17029; X_Im[501]=32'd15716; X_Im[1013]=32'd5513; X_Im[13]=32'd6176; X_Im[525]=32'd8068; X_Im[269]=-32'd17029; X_Im[781]=-32'd2672; X_Im[141]=-32'd1375; X_Im[653]=-32'd5924; X_Im[397]=-32'd4235; X_Im[909]=-32'd1369; X_Im[77]=-32'd372; X_Im[589]=32'd1316; X_Im[333]=32'd2306; X_Im[845]=32'd12769; X_Im[205]=32'd4959; X_Im[717]=32'd7091; X_Im[461]=32'd6966; X_Im[973]=32'd4202; X_Im[45]=32'd2408; X_Im[557]=32'd7040; X_Im[301]=-32'd3541; X_Im[813]=32'd3416; X_Im[173]=-32'd412; X_Im[685]=-32'd2085; X_Im[429]=-32'd21317; X_Im[941]=-32'd1411; X_Im[109]=32'd39175; X_Im[621]=32'd11007; X_Im[365]=32'd6800; X_Im[877]=-32'd3262; X_Im[237]=32'd10580; X_Im[749]=32'd2488; X_Im[493]=32'd13702; X_Im[1005]=32'd9133; X_Im[29]=32'd9143; X_Im[541]=32'd4612; X_Im[285]=32'd5407; X_Im[797]=32'd15490; X_Im[157]=-32'd2578; X_Im[669]=32'd29632; X_Im[413]=-32'd22921; X_Im[925]=32'd23781; X_Im[93]=32'd14740; X_Im[605]=32'd1199; X_Im[349]=-32'd4875; X_Im[861]=-32'd10964; X_Im[221]=32'd857; X_Im[733]=-32'd2246; X_Im[477]=-32'd5730; X_Im[989]=32'd10534; X_Im[61]=32'd11436; X_Im[573]=32'd13946; X_Im[317]=32'd39729; X_Im[829]=-32'd67060; X_Im[189]=32'd21451; X_Im[701]=-32'd19877; X_Im[445]=-32'd8936; X_Im[957]=-32'd16399; X_Im[125]=32'd5325; X_Im[637]=32'd12687; X_Im[381]=32'd7979; X_Im[893]=32'd1942; X_Im[253]=-32'd1441; X_Im[765]=32'd7941; X_Im[509]=-32'd4283; X_Im[1021]=-32'd658; X_Im[3]=32'd2824; X_Im[515]=-32'd7721; X_Im[259]=-32'd5393; X_Im[771]=32'd3797; X_Im[131]=-32'd3903; X_Im[643]=32'd2923; X_Im[387]=32'd2390; X_Im[899]=32'd4159; X_Im[67]=32'd1652; X_Im[579]=-32'd93; X_Im[323]=32'd6068; X_Im[835]=32'd4814; X_Im[195]=32'd2579; X_Im[707]=-32'd543; X_Im[451]=-32'd15040; X_Im[963]=32'd3686; X_Im[35]=32'd5725; X_Im[547]=32'd7724; X_Im[291]=32'd5439; X_Im[803]=32'd16467; X_Im[163]=-32'd2644; X_Im[675]=32'd15006; X_Im[419]=32'd3671; X_Im[931]=32'd11132; X_Im[99]=32'd4480; X_Im[611]=32'd1958; X_Im[355]=32'd647; X_Im[867]=-32'd759; X_Im[227]=32'd1380; X_Im[739]=32'd4288; X_Im[483]=32'd7358; X_Im[995]=32'd7961; X_Im[19]=32'd1015; X_Im[531]=32'd11491; X_Im[275]=-32'd9592; X_Im[787]=32'd6244; X_Im[147]=32'd5421; X_Im[659]=32'd10742; X_Im[403]=32'd12617; X_Im[915]=32'd13536; X_Im[83]=32'd7149; X_Im[595]=32'd12952; X_Im[339]=32'd11902; X_Im[851]=32'd18114; X_Im[211]=-32'd1116; X_Im[723]=32'd11523; X_Im[467]=32'd10890; X_Im[979]=32'd11450; X_Im[51]=32'd13366; X_Im[563]=32'd19440; X_Im[307]=32'd20123; X_Im[819]=32'd13828; X_Im[179]=32'd25585; X_Im[691]=32'd37908; X_Im[435]=-32'd4902; X_Im[947]=32'd134452; X_Im[115]=-32'd58461; X_Im[627]=-32'd63798; X_Im[371]=-32'd98891; X_Im[883]=-32'd64467; X_Im[243]=-32'd30560; X_Im[755]=-32'd22139; X_Im[499]=-32'd12192; X_Im[1011]=-32'd16888; X_Im[11]=-32'd1345; X_Im[523]=-32'd10858; X_Im[267]=-32'd4871; X_Im[779]=32'd15558; X_Im[139]=-32'd11756; X_Im[651]=-32'd25003; X_Im[395]=-32'd2570; X_Im[907]=32'd1846; X_Im[75]=-32'd11040; X_Im[587]=-32'd1474; X_Im[331]=32'd2780; X_Im[843]=-32'd1537; X_Im[203]=-32'd13251; X_Im[715]=-32'd19053; X_Im[459]=32'd17162; X_Im[971]=-32'd10031; X_Im[43]=-32'd2011; X_Im[555]=-32'd686; X_Im[299]=32'd1992; X_Im[811]=-32'd6524; X_Im[171]=-32'd5402; X_Im[683]=32'd3625; X_Im[427]=-32'd8437; X_Im[939]=32'd3376; X_Im[107]=-32'd7049; X_Im[619]=-32'd5613; X_Im[363]=-32'd9738; X_Im[875]=-32'd8129; X_Im[235]=-32'd14901; X_Im[747]=-32'd3204; X_Im[491]=-32'd10007; X_Im[1003]=32'd45472; X_Im[27]=32'd30401; X_Im[539]=-32'd73732; X_Im[283]=32'd38556; X_Im[795]=32'd25667; X_Im[155]=32'd4537; X_Im[667]=32'd676; X_Im[411]=32'd89; X_Im[923]=-32'd5153; X_Im[91]=32'd2636; X_Im[603]=-32'd4257; X_Im[347]=-32'd3011; X_Im[859]=-32'd766; X_Im[219]=32'd339; X_Im[731]=32'd1974; X_Im[475]=-32'd1; X_Im[987]=-32'd1260; X_Im[59]=32'd5964; X_Im[571]=-32'd7477; X_Im[315]=-32'd10751; X_Im[827]=-32'd42849; X_Im[187]=-32'd17405; X_Im[699]=-32'd9077; X_Im[443]=-32'd5862; X_Im[955]=-32'd13203; X_Im[123]=32'd17815; X_Im[635]=-32'd148481; X_Im[379]=32'd175459; X_Im[891]=32'd29326; X_Im[251]=-32'd77885; X_Im[763]=-32'd43848; X_Im[507]=-32'd24502; X_Im[1019]=-32'd18947; X_Im[7]=-32'd14000; X_Im[519]=-32'd16925; X_Im[263]=-32'd17927; X_Im[775]=-32'd22138; X_Im[135]=-32'd21897; X_Im[647]=-32'd8339; X_Im[391]=-32'd32457; X_Im[903]=-32'd4768; X_Im[71]=-32'd159144; X_Im[583]=-32'd133139; X_Im[327]=32'd30338; X_Im[839]=32'd114821; X_Im[199]=32'd54085; X_Im[711]=32'd32225; X_Im[455]=32'd32568; X_Im[967]=32'd15082; X_Im[39]=32'd32539; X_Im[551]=32'd2572; X_Im[295]=32'd8343; X_Im[807]=32'd5188; X_Im[167]=-32'd4870; X_Im[679]=-32'd8519; X_Im[423]=-32'd22830; X_Im[935]=32'd11776; X_Im[103]=32'd21730; X_Im[615]=32'd5380; X_Im[359]=32'd8961; X_Im[871]=32'd991; X_Im[231]=-32'd2601; X_Im[743]=32'd1126; X_Im[487]=-32'd6873; X_Im[999]=32'd1057; X_Im[23]=32'd11538; X_Im[535]=32'd1563; X_Im[279]=32'd25124; X_Im[791]=32'd7105; X_Im[151]=32'd24689; X_Im[663]=32'd30190; X_Im[407]=32'd34823; X_Im[919]=-32'd66525; X_Im[87]=-32'd46374; X_Im[599]=-32'd11844; X_Im[343]=-32'd9496; X_Im[855]=-32'd14039; X_Im[215]=-32'd12639; X_Im[727]=-32'd23195; X_Im[471]=-32'd34833; X_Im[983]=-32'd75688; X_Im[55]=-32'd70691; X_Im[567]=32'd183414; X_Im[311]=32'd64712; X_Im[823]=32'd40605; X_Im[183]=32'd27931; X_Im[695]=32'd33190; X_Im[439]=32'd22629; X_Im[951]=32'd10093; X_Im[119]=32'd55297; X_Im[631]=32'd63305; X_Im[375]=-32'd1668; X_Im[887]=-32'd4696; X_Im[247]=-32'd151433; X_Im[759]=32'd714901; X_Im[503]=-32'd124522; X_Im[1015]=-32'd6967; X_Im[15]=32'd10776; X_Im[527]=-32'd4488; X_Im[271]=-32'd8026; X_Im[783]=32'd5077; X_Im[143]=-32'd6643; X_Im[655]=32'd182053; X_Im[399]=32'd88372; X_Im[911]=32'd4368; X_Im[79]=32'd44533; X_Im[591]=32'd34272; X_Im[335]=32'd32459; X_Im[847]=-32'd87188; X_Im[207]=-32'd11192; X_Im[719]=32'd22785; X_Im[463]=32'd7730; X_Im[975]=32'd30607; X_Im[47]=32'd26484; X_Im[559]=-32'd85512; X_Im[303]=32'd5987; X_Im[815]=-32'd40748; X_Im[175]=32'd22530; X_Im[687]=32'd66258; X_Im[431]=32'd77472; X_Im[943]=32'd114939; X_Im[111]=32'd332002; X_Im[623]=-32'd611736; X_Im[367]=-32'd154365; X_Im[879]=-32'd87548; X_Im[239]=-32'd67934; X_Im[751]=-32'd88522; X_Im[495]=-32'd52457; X_Im[1007]=-32'd46075; X_Im[31]=-32'd37022; X_Im[543]=-32'd36200; X_Im[287]=-32'd31296; X_Im[799]=-32'd25853; X_Im[159]=-32'd28244; X_Im[671]=-32'd20701; X_Im[415]=32'd11679; X_Im[927]=-32'd8041; X_Im[95]=-32'd12985; X_Im[607]=32'd17590; X_Im[351]=-32'd21141; X_Im[863]=-32'd19111; X_Im[223]=-32'd46940; X_Im[735]=-32'd42162; X_Im[479]=-32'd64934; X_Im[991]=-32'd4976; X_Im[63]=-32'd6583; X_Im[575]=-32'd15022; X_Im[319]=32'd12300; X_Im[831]=-32'd94271; X_Im[191]=-32'd25657; X_Im[703]=-32'd12968; X_Im[447]=-32'd35545; X_Im[959]=-32'd139265; X_Im[127]=32'd40194; X_Im[639]=-32'd48603; X_Im[383]=32'd73376; X_Im[895]=32'd34136; X_Im[255]=32'd30790; X_Im[767]=32'd28663; X_Im[511]=32'd12913; X_Im[1023]=32'd1486;
		#10
		Reset = 0;
		#10
		
		Start = 1;
		#130
		Start = 0;
	end

endmodule