`timescale 1ns / 1ps

module FFT1024_tb_v;
	parameter PRE = 32;
		
	reg Clk;
	reg Reset, Start, Ack;
	reg signed [PRE-1:0] X_Re [1023:0];
	reg signed [PRE-1:0] X_Im [1023:0];
	
	// Outputs
	wire [PRE*1024-1:0] Y_Re_out;
	wire [PRE*1024-1:0] Y_Im_out;
	wire [3:0] state;
	wire Done;
	
	// Internal
	wire [32*1024-1:0] X_Re_Packed = { X_Re[1023], X_Re[1022], X_Re[1021], X_Re[1020], X_Re[1019], X_Re[1018], X_Re[1017], X_Re[1016], X_Re[1015], X_Re[1014], X_Re[1013], X_Re[1012], X_Re[1011], X_Re[1010], X_Re[1009], X_Re[1008], X_Re[1007], X_Re[1006], X_Re[1005], X_Re[1004], X_Re[1003], X_Re[1002], X_Re[1001], X_Re[1000], X_Re[999], X_Re[998], X_Re[997], X_Re[996], X_Re[995], X_Re[994], X_Re[993], X_Re[992], X_Re[991], X_Re[990], X_Re[989], X_Re[988], X_Re[987], X_Re[986], X_Re[985], X_Re[984], X_Re[983], X_Re[982], X_Re[981], X_Re[980], X_Re[979], X_Re[978], X_Re[977], X_Re[976], X_Re[975], X_Re[974], X_Re[973], X_Re[972], X_Re[971], X_Re[970], X_Re[969], X_Re[968], X_Re[967], X_Re[966], X_Re[965], X_Re[964], X_Re[963], X_Re[962], X_Re[961], X_Re[960], X_Re[959], X_Re[958], X_Re[957], X_Re[956], X_Re[955], X_Re[954], X_Re[953], X_Re[952], X_Re[951], X_Re[950], X_Re[949], X_Re[948], X_Re[947], X_Re[946], X_Re[945], X_Re[944], X_Re[943], X_Re[942], X_Re[941], X_Re[940], X_Re[939], X_Re[938], X_Re[937], X_Re[936], X_Re[935], X_Re[934], X_Re[933], X_Re[932], X_Re[931], X_Re[930], X_Re[929], X_Re[928], X_Re[927], X_Re[926], X_Re[925], X_Re[924], X_Re[923], X_Re[922], X_Re[921], X_Re[920], X_Re[919], X_Re[918], X_Re[917], X_Re[916], X_Re[915], X_Re[914], X_Re[913], X_Re[912], X_Re[911], X_Re[910], X_Re[909], X_Re[908], X_Re[907], X_Re[906], X_Re[905], X_Re[904], X_Re[903], X_Re[902], X_Re[901], X_Re[900], X_Re[899], X_Re[898], X_Re[897], X_Re[896], X_Re[895], X_Re[894], X_Re[893], X_Re[892], X_Re[891], X_Re[890], X_Re[889], X_Re[888], X_Re[887], X_Re[886], X_Re[885], X_Re[884], X_Re[883], X_Re[882], X_Re[881], X_Re[880], X_Re[879], X_Re[878], X_Re[877], X_Re[876], X_Re[875], X_Re[874], X_Re[873], X_Re[872], X_Re[871], X_Re[870], X_Re[869], X_Re[868], X_Re[867], X_Re[866], X_Re[865], X_Re[864], X_Re[863], X_Re[862], X_Re[861], X_Re[860], X_Re[859], X_Re[858], X_Re[857], X_Re[856], X_Re[855], X_Re[854], X_Re[853], X_Re[852], X_Re[851], X_Re[850], X_Re[849], X_Re[848], X_Re[847], X_Re[846], X_Re[845], X_Re[844], X_Re[843], X_Re[842], X_Re[841], X_Re[840], X_Re[839], X_Re[838], X_Re[837], X_Re[836], X_Re[835], X_Re[834], X_Re[833], X_Re[832], X_Re[831], X_Re[830], X_Re[829], X_Re[828], X_Re[827], X_Re[826], X_Re[825], X_Re[824], X_Re[823], X_Re[822], X_Re[821], X_Re[820], X_Re[819], X_Re[818], X_Re[817], X_Re[816], X_Re[815], X_Re[814], X_Re[813], X_Re[812], X_Re[811], X_Re[810], X_Re[809], X_Re[808], X_Re[807], X_Re[806], X_Re[805], X_Re[804], X_Re[803], X_Re[802], X_Re[801], X_Re[800], X_Re[799], X_Re[798], X_Re[797], X_Re[796], X_Re[795], X_Re[794], X_Re[793], X_Re[792], X_Re[791], X_Re[790], X_Re[789], X_Re[788], X_Re[787], X_Re[786], X_Re[785], X_Re[784], X_Re[783], X_Re[782], X_Re[781], X_Re[780], X_Re[779], X_Re[778], X_Re[777], X_Re[776], X_Re[775], X_Re[774], X_Re[773], X_Re[772], X_Re[771], X_Re[770], X_Re[769], X_Re[768], X_Re[767], X_Re[766], X_Re[765], X_Re[764], X_Re[763], X_Re[762], X_Re[761], X_Re[760], X_Re[759], X_Re[758], X_Re[757], X_Re[756], X_Re[755], X_Re[754], X_Re[753], X_Re[752], X_Re[751], X_Re[750], X_Re[749], X_Re[748], X_Re[747], X_Re[746], X_Re[745], X_Re[744], X_Re[743], X_Re[742], X_Re[741], X_Re[740], X_Re[739], X_Re[738], X_Re[737], X_Re[736], X_Re[735], X_Re[734], X_Re[733], X_Re[732], X_Re[731], X_Re[730], X_Re[729], X_Re[728], X_Re[727], X_Re[726], X_Re[725], X_Re[724], X_Re[723], X_Re[722], X_Re[721], X_Re[720], X_Re[719], X_Re[718], X_Re[717], X_Re[716], X_Re[715], X_Re[714], X_Re[713], X_Re[712], X_Re[711], X_Re[710], X_Re[709], X_Re[708], X_Re[707], X_Re[706], X_Re[705], X_Re[704], X_Re[703], X_Re[702], X_Re[701], X_Re[700], X_Re[699], X_Re[698], X_Re[697], X_Re[696], X_Re[695], X_Re[694], X_Re[693], X_Re[692], X_Re[691], X_Re[690], X_Re[689], X_Re[688], X_Re[687], X_Re[686], X_Re[685], X_Re[684], X_Re[683], X_Re[682], X_Re[681], X_Re[680], X_Re[679], X_Re[678], X_Re[677], X_Re[676], X_Re[675], X_Re[674], X_Re[673], X_Re[672], X_Re[671], X_Re[670], X_Re[669], X_Re[668], X_Re[667], X_Re[666], X_Re[665], X_Re[664], X_Re[663], X_Re[662], X_Re[661], X_Re[660], X_Re[659], X_Re[658], X_Re[657], X_Re[656], X_Re[655], X_Re[654], X_Re[653], X_Re[652], X_Re[651], X_Re[650], X_Re[649], X_Re[648], X_Re[647], X_Re[646], X_Re[645], X_Re[644], X_Re[643], X_Re[642], X_Re[641], X_Re[640], X_Re[639], X_Re[638], X_Re[637], X_Re[636], X_Re[635], X_Re[634], X_Re[633], X_Re[632], X_Re[631], X_Re[630], X_Re[629], X_Re[628], X_Re[627], X_Re[626], X_Re[625], X_Re[624], X_Re[623], X_Re[622], X_Re[621], X_Re[620], X_Re[619], X_Re[618], X_Re[617], X_Re[616], X_Re[615], X_Re[614], X_Re[613], X_Re[612], X_Re[611], X_Re[610], X_Re[609], X_Re[608], X_Re[607], X_Re[606], X_Re[605], X_Re[604], X_Re[603], X_Re[602], X_Re[601], X_Re[600], X_Re[599], X_Re[598], X_Re[597], X_Re[596], X_Re[595], X_Re[594], X_Re[593], X_Re[592], X_Re[591], X_Re[590], X_Re[589], X_Re[588], X_Re[587], X_Re[586], X_Re[585], X_Re[584], X_Re[583], X_Re[582], X_Re[581], X_Re[580], X_Re[579], X_Re[578], X_Re[577], X_Re[576], X_Re[575], X_Re[574], X_Re[573], X_Re[572], X_Re[571], X_Re[570], X_Re[569], X_Re[568], X_Re[567], X_Re[566], X_Re[565], X_Re[564], X_Re[563], X_Re[562], X_Re[561], X_Re[560], X_Re[559], X_Re[558], X_Re[557], X_Re[556], X_Re[555], X_Re[554], X_Re[553], X_Re[552], X_Re[551], X_Re[550], X_Re[549], X_Re[548], X_Re[547], X_Re[546], X_Re[545], X_Re[544], X_Re[543], X_Re[542], X_Re[541], X_Re[540], X_Re[539], X_Re[538], X_Re[537], X_Re[536], X_Re[535], X_Re[534], X_Re[533], X_Re[532], X_Re[531], X_Re[530], X_Re[529], X_Re[528], X_Re[527], X_Re[526], X_Re[525], X_Re[524], X_Re[523], X_Re[522], X_Re[521], X_Re[520], X_Re[519], X_Re[518], X_Re[517], X_Re[516], X_Re[515], X_Re[514], X_Re[513], X_Re[512], X_Re[511], X_Re[510], X_Re[509], X_Re[508], X_Re[507], X_Re[506], X_Re[505], X_Re[504], X_Re[503], X_Re[502], X_Re[501], X_Re[500], X_Re[499], X_Re[498], X_Re[497], X_Re[496], X_Re[495], X_Re[494], X_Re[493], X_Re[492], X_Re[491], X_Re[490], X_Re[489], X_Re[488], X_Re[487], X_Re[486], X_Re[485], X_Re[484], X_Re[483], X_Re[482], X_Re[481], X_Re[480], X_Re[479], X_Re[478], X_Re[477], X_Re[476], X_Re[475], X_Re[474], X_Re[473], X_Re[472], X_Re[471], X_Re[470], X_Re[469], X_Re[468], X_Re[467], X_Re[466], X_Re[465], X_Re[464], X_Re[463], X_Re[462], X_Re[461], X_Re[460], X_Re[459], X_Re[458], X_Re[457], X_Re[456], X_Re[455], X_Re[454], X_Re[453], X_Re[452], X_Re[451], X_Re[450], X_Re[449], X_Re[448], X_Re[447], X_Re[446], X_Re[445], X_Re[444], X_Re[443], X_Re[442], X_Re[441], X_Re[440], X_Re[439], X_Re[438], X_Re[437], X_Re[436], X_Re[435], X_Re[434], X_Re[433], X_Re[432], X_Re[431], X_Re[430], X_Re[429], X_Re[428], X_Re[427], X_Re[426], X_Re[425], X_Re[424], X_Re[423], X_Re[422], X_Re[421], X_Re[420], X_Re[419], X_Re[418], X_Re[417], X_Re[416], X_Re[415], X_Re[414], X_Re[413], X_Re[412], X_Re[411], X_Re[410], X_Re[409], X_Re[408], X_Re[407], X_Re[406], X_Re[405], X_Re[404], X_Re[403], X_Re[402], X_Re[401], X_Re[400], X_Re[399], X_Re[398], X_Re[397], X_Re[396], X_Re[395], X_Re[394], X_Re[393], X_Re[392], X_Re[391], X_Re[390], X_Re[389], X_Re[388], X_Re[387], X_Re[386], X_Re[385], X_Re[384], X_Re[383], X_Re[382], X_Re[381], X_Re[380], X_Re[379], X_Re[378], X_Re[377], X_Re[376], X_Re[375], X_Re[374], X_Re[373], X_Re[372], X_Re[371], X_Re[370], X_Re[369], X_Re[368], X_Re[367], X_Re[366], X_Re[365], X_Re[364], X_Re[363], X_Re[362], X_Re[361], X_Re[360], X_Re[359], X_Re[358], X_Re[357], X_Re[356], X_Re[355], X_Re[354], X_Re[353], X_Re[352], X_Re[351], X_Re[350], X_Re[349], X_Re[348], X_Re[347], X_Re[346], X_Re[345], X_Re[344], X_Re[343], X_Re[342], X_Re[341], X_Re[340], X_Re[339], X_Re[338], X_Re[337], X_Re[336], X_Re[335], X_Re[334], X_Re[333], X_Re[332], X_Re[331], X_Re[330], X_Re[329], X_Re[328], X_Re[327], X_Re[326], X_Re[325], X_Re[324], X_Re[323], X_Re[322], X_Re[321], X_Re[320], X_Re[319], X_Re[318], X_Re[317], X_Re[316], X_Re[315], X_Re[314], X_Re[313], X_Re[312], X_Re[311], X_Re[310], X_Re[309], X_Re[308], X_Re[307], X_Re[306], X_Re[305], X_Re[304], X_Re[303], X_Re[302], X_Re[301], X_Re[300], X_Re[299], X_Re[298], X_Re[297], X_Re[296], X_Re[295], X_Re[294], X_Re[293], X_Re[292], X_Re[291], X_Re[290], X_Re[289], X_Re[288], X_Re[287], X_Re[286], X_Re[285], X_Re[284], X_Re[283], X_Re[282], X_Re[281], X_Re[280], X_Re[279], X_Re[278], X_Re[277], X_Re[276], X_Re[275], X_Re[274], X_Re[273], X_Re[272], X_Re[271], X_Re[270], X_Re[269], X_Re[268], X_Re[267], X_Re[266], X_Re[265], X_Re[264], X_Re[263], X_Re[262], X_Re[261], X_Re[260], X_Re[259], X_Re[258], X_Re[257], X_Re[256], X_Re[255], X_Re[254], X_Re[253], X_Re[252], X_Re[251], X_Re[250], X_Re[249], X_Re[248], X_Re[247], X_Re[246], X_Re[245], X_Re[244], X_Re[243], X_Re[242], X_Re[241], X_Re[240], X_Re[239], X_Re[238], X_Re[237], X_Re[236], X_Re[235], X_Re[234], X_Re[233], X_Re[232], X_Re[231], X_Re[230], X_Re[229], X_Re[228], X_Re[227], X_Re[226], X_Re[225], X_Re[224], X_Re[223], X_Re[222], X_Re[221], X_Re[220], X_Re[219], X_Re[218], X_Re[217], X_Re[216], X_Re[215], X_Re[214], X_Re[213], X_Re[212], X_Re[211], X_Re[210], X_Re[209], X_Re[208], X_Re[207], X_Re[206], X_Re[205], X_Re[204], X_Re[203], X_Re[202], X_Re[201], X_Re[200], X_Re[199], X_Re[198], X_Re[197], X_Re[196], X_Re[195], X_Re[194], X_Re[193], X_Re[192], X_Re[191], X_Re[190], X_Re[189], X_Re[188], X_Re[187], X_Re[186], X_Re[185], X_Re[184], X_Re[183], X_Re[182], X_Re[181], X_Re[180], X_Re[179], X_Re[178], X_Re[177], X_Re[176], X_Re[175], X_Re[174], X_Re[173], X_Re[172], X_Re[171], X_Re[170], X_Re[169], X_Re[168], X_Re[167], X_Re[166], X_Re[165], X_Re[164], X_Re[163], X_Re[162], X_Re[161], X_Re[160], X_Re[159], X_Re[158], X_Re[157], X_Re[156], X_Re[155], X_Re[154], X_Re[153], X_Re[152], X_Re[151], X_Re[150], X_Re[149], X_Re[148], X_Re[147], X_Re[146], X_Re[145], X_Re[144], X_Re[143], X_Re[142], X_Re[141], X_Re[140], X_Re[139], X_Re[138], X_Re[137], X_Re[136], X_Re[135], X_Re[134], X_Re[133], X_Re[132], X_Re[131], X_Re[130], X_Re[129], X_Re[128], X_Re[127], X_Re[126], X_Re[125], X_Re[124], X_Re[123], X_Re[122], X_Re[121], X_Re[120], X_Re[119], X_Re[118], X_Re[117], X_Re[116], X_Re[115], X_Re[114], X_Re[113], X_Re[112], X_Re[111], X_Re[110], X_Re[109], X_Re[108], X_Re[107], X_Re[106], X_Re[105], X_Re[104], X_Re[103], X_Re[102], X_Re[101], X_Re[100], X_Re[99], X_Re[98], X_Re[97], X_Re[96], X_Re[95], X_Re[94], X_Re[93], X_Re[92], X_Re[91], X_Re[90], X_Re[89], X_Re[88], X_Re[87], X_Re[86], X_Re[85], X_Re[84], X_Re[83], X_Re[82], X_Re[81], X_Re[80], X_Re[79], X_Re[78], X_Re[77], X_Re[76], X_Re[75], X_Re[74], X_Re[73], X_Re[72], X_Re[71], X_Re[70], X_Re[69], X_Re[68], X_Re[67], X_Re[66], X_Re[65], X_Re[64], X_Re[63], X_Re[62], X_Re[61], X_Re[60], X_Re[59], X_Re[58], X_Re[57], X_Re[56], X_Re[55], X_Re[54], X_Re[53], X_Re[52], X_Re[51], X_Re[50], X_Re[49], X_Re[48], X_Re[47], X_Re[46], X_Re[45], X_Re[44], X_Re[43], X_Re[42], X_Re[41], X_Re[40], X_Re[39], X_Re[38], X_Re[37], X_Re[36], X_Re[35], X_Re[34], X_Re[33], X_Re[32], X_Re[31], X_Re[30], X_Re[29], X_Re[28], X_Re[27], X_Re[26], X_Re[25], X_Re[24], X_Re[23], X_Re[22], X_Re[21], X_Re[20], X_Re[19], X_Re[18], X_Re[17], X_Re[16], X_Re[15], X_Re[14], X_Re[13], X_Re[12], X_Re[11], X_Re[10], X_Re[9], X_Re[8], X_Re[7], X_Re[6], X_Re[5], X_Re[4], X_Re[3], X_Re[2], X_Re[1], X_Re[0]};
	wire [1024*16-1:0] X_Im_Packed = { X_Im[1023], X_Im[1022], X_Im[1021], X_Im[1020], X_Im[1019], X_Im[1018], X_Im[1017], X_Im[1016], X_Im[1015], X_Im[1014], X_Im[1013], X_Im[1012], X_Im[1011], X_Im[1010], X_Im[1009], X_Im[1008], X_Im[1007], X_Im[1006], X_Im[1005], X_Im[1004], X_Im[1003], X_Im[1002], X_Im[1001], X_Im[1000], X_Im[999], X_Im[998], X_Im[997], X_Im[996], X_Im[995], X_Im[994], X_Im[993], X_Im[992], X_Im[991], X_Im[990], X_Im[989], X_Im[988], X_Im[987], X_Im[986], X_Im[985], X_Im[984], X_Im[983], X_Im[982], X_Im[981], X_Im[980], X_Im[979], X_Im[978], X_Im[977], X_Im[976], X_Im[975], X_Im[974], X_Im[973], X_Im[972], X_Im[971], X_Im[970], X_Im[969], X_Im[968], X_Im[967], X_Im[966], X_Im[965], X_Im[964], X_Im[963], X_Im[962], X_Im[961], X_Im[960], X_Im[959], X_Im[958], X_Im[957], X_Im[956], X_Im[955], X_Im[954], X_Im[953], X_Im[952], X_Im[951], X_Im[950], X_Im[949], X_Im[948], X_Im[947], X_Im[946], X_Im[945], X_Im[944], X_Im[943], X_Im[942], X_Im[941], X_Im[940], X_Im[939], X_Im[938], X_Im[937], X_Im[936], X_Im[935], X_Im[934], X_Im[933], X_Im[932], X_Im[931], X_Im[930], X_Im[929], X_Im[928], X_Im[927], X_Im[926], X_Im[925], X_Im[924], X_Im[923], X_Im[922], X_Im[921], X_Im[920], X_Im[919], X_Im[918], X_Im[917], X_Im[916], X_Im[915], X_Im[914], X_Im[913], X_Im[912], X_Im[911], X_Im[910], X_Im[909], X_Im[908], X_Im[907], X_Im[906], X_Im[905], X_Im[904], X_Im[903], X_Im[902], X_Im[901], X_Im[900], X_Im[899], X_Im[898], X_Im[897], X_Im[896], X_Im[895], X_Im[894], X_Im[893], X_Im[892], X_Im[891], X_Im[890], X_Im[889], X_Im[888], X_Im[887], X_Im[886], X_Im[885], X_Im[884], X_Im[883], X_Im[882], X_Im[881], X_Im[880], X_Im[879], X_Im[878], X_Im[877], X_Im[876], X_Im[875], X_Im[874], X_Im[873], X_Im[872], X_Im[871], X_Im[870], X_Im[869], X_Im[868], X_Im[867], X_Im[866], X_Im[865], X_Im[864], X_Im[863], X_Im[862], X_Im[861], X_Im[860], X_Im[859], X_Im[858], X_Im[857], X_Im[856], X_Im[855], X_Im[854], X_Im[853], X_Im[852], X_Im[851], X_Im[850], X_Im[849], X_Im[848], X_Im[847], X_Im[846], X_Im[845], X_Im[844], X_Im[843], X_Im[842], X_Im[841], X_Im[840], X_Im[839], X_Im[838], X_Im[837], X_Im[836], X_Im[835], X_Im[834], X_Im[833], X_Im[832], X_Im[831], X_Im[830], X_Im[829], X_Im[828], X_Im[827], X_Im[826], X_Im[825], X_Im[824], X_Im[823], X_Im[822], X_Im[821], X_Im[820], X_Im[819], X_Im[818], X_Im[817], X_Im[816], X_Im[815], X_Im[814], X_Im[813], X_Im[812], X_Im[811], X_Im[810], X_Im[809], X_Im[808], X_Im[807], X_Im[806], X_Im[805], X_Im[804], X_Im[803], X_Im[802], X_Im[801], X_Im[800], X_Im[799], X_Im[798], X_Im[797], X_Im[796], X_Im[795], X_Im[794], X_Im[793], X_Im[792], X_Im[791], X_Im[790], X_Im[789], X_Im[788], X_Im[787], X_Im[786], X_Im[785], X_Im[784], X_Im[783], X_Im[782], X_Im[781], X_Im[780], X_Im[779], X_Im[778], X_Im[777], X_Im[776], X_Im[775], X_Im[774], X_Im[773], X_Im[772], X_Im[771], X_Im[770], X_Im[769], X_Im[768], X_Im[767], X_Im[766], X_Im[765], X_Im[764], X_Im[763], X_Im[762], X_Im[761], X_Im[760], X_Im[759], X_Im[758], X_Im[757], X_Im[756], X_Im[755], X_Im[754], X_Im[753], X_Im[752], X_Im[751], X_Im[750], X_Im[749], X_Im[748], X_Im[747], X_Im[746], X_Im[745], X_Im[744], X_Im[743], X_Im[742], X_Im[741], X_Im[740], X_Im[739], X_Im[738], X_Im[737], X_Im[736], X_Im[735], X_Im[734], X_Im[733], X_Im[732], X_Im[731], X_Im[730], X_Im[729], X_Im[728], X_Im[727], X_Im[726], X_Im[725], X_Im[724], X_Im[723], X_Im[722], X_Im[721], X_Im[720], X_Im[719], X_Im[718], X_Im[717], X_Im[716], X_Im[715], X_Im[714], X_Im[713], X_Im[712], X_Im[711], X_Im[710], X_Im[709], X_Im[708], X_Im[707], X_Im[706], X_Im[705], X_Im[704], X_Im[703], X_Im[702], X_Im[701], X_Im[700], X_Im[699], X_Im[698], X_Im[697], X_Im[696], X_Im[695], X_Im[694], X_Im[693], X_Im[692], X_Im[691], X_Im[690], X_Im[689], X_Im[688], X_Im[687], X_Im[686], X_Im[685], X_Im[684], X_Im[683], X_Im[682], X_Im[681], X_Im[680], X_Im[679], X_Im[678], X_Im[677], X_Im[676], X_Im[675], X_Im[674], X_Im[673], X_Im[672], X_Im[671], X_Im[670], X_Im[669], X_Im[668], X_Im[667], X_Im[666], X_Im[665], X_Im[664], X_Im[663], X_Im[662], X_Im[661], X_Im[660], X_Im[659], X_Im[658], X_Im[657], X_Im[656], X_Im[655], X_Im[654], X_Im[653], X_Im[652], X_Im[651], X_Im[650], X_Im[649], X_Im[648], X_Im[647], X_Im[646], X_Im[645], X_Im[644], X_Im[643], X_Im[642], X_Im[641], X_Im[640], X_Im[639], X_Im[638], X_Im[637], X_Im[636], X_Im[635], X_Im[634], X_Im[633], X_Im[632], X_Im[631], X_Im[630], X_Im[629], X_Im[628], X_Im[627], X_Im[626], X_Im[625], X_Im[624], X_Im[623], X_Im[622], X_Im[621], X_Im[620], X_Im[619], X_Im[618], X_Im[617], X_Im[616], X_Im[615], X_Im[614], X_Im[613], X_Im[612], X_Im[611], X_Im[610], X_Im[609], X_Im[608], X_Im[607], X_Im[606], X_Im[605], X_Im[604], X_Im[603], X_Im[602], X_Im[601], X_Im[600], X_Im[599], X_Im[598], X_Im[597], X_Im[596], X_Im[595], X_Im[594], X_Im[593], X_Im[592], X_Im[591], X_Im[590], X_Im[589], X_Im[588], X_Im[587], X_Im[586], X_Im[585], X_Im[584], X_Im[583], X_Im[582], X_Im[581], X_Im[580], X_Im[579], X_Im[578], X_Im[577], X_Im[576], X_Im[575], X_Im[574], X_Im[573], X_Im[572], X_Im[571], X_Im[570], X_Im[569], X_Im[568], X_Im[567], X_Im[566], X_Im[565], X_Im[564], X_Im[563], X_Im[562], X_Im[561], X_Im[560], X_Im[559], X_Im[558], X_Im[557], X_Im[556], X_Im[555], X_Im[554], X_Im[553], X_Im[552], X_Im[551], X_Im[550], X_Im[549], X_Im[548], X_Im[547], X_Im[546], X_Im[545], X_Im[544], X_Im[543], X_Im[542], X_Im[541], X_Im[540], X_Im[539], X_Im[538], X_Im[537], X_Im[536], X_Im[535], X_Im[534], X_Im[533], X_Im[532], X_Im[531], X_Im[530], X_Im[529], X_Im[528], X_Im[527], X_Im[526], X_Im[525], X_Im[524], X_Im[523], X_Im[522], X_Im[521], X_Im[520], X_Im[519], X_Im[518], X_Im[517], X_Im[516], X_Im[515], X_Im[514], X_Im[513], X_Im[512], X_Im[511], X_Im[510], X_Im[509], X_Im[508], X_Im[507], X_Im[506], X_Im[505], X_Im[504], X_Im[503], X_Im[502], X_Im[501], X_Im[500], X_Im[499], X_Im[498], X_Im[497], X_Im[496], X_Im[495], X_Im[494], X_Im[493], X_Im[492], X_Im[491], X_Im[490], X_Im[489], X_Im[488], X_Im[487], X_Im[486], X_Im[485], X_Im[484], X_Im[483], X_Im[482], X_Im[481], X_Im[480], X_Im[479], X_Im[478], X_Im[477], X_Im[476], X_Im[475], X_Im[474], X_Im[473], X_Im[472], X_Im[471], X_Im[470], X_Im[469], X_Im[468], X_Im[467], X_Im[466], X_Im[465], X_Im[464], X_Im[463], X_Im[462], X_Im[461], X_Im[460], X_Im[459], X_Im[458], X_Im[457], X_Im[456], X_Im[455], X_Im[454], X_Im[453], X_Im[452], X_Im[451], X_Im[450], X_Im[449], X_Im[448], X_Im[447], X_Im[446], X_Im[445], X_Im[444], X_Im[443], X_Im[442], X_Im[441], X_Im[440], X_Im[439], X_Im[438], X_Im[437], X_Im[436], X_Im[435], X_Im[434], X_Im[433], X_Im[432], X_Im[431], X_Im[430], X_Im[429], X_Im[428], X_Im[427], X_Im[426], X_Im[425], X_Im[424], X_Im[423], X_Im[422], X_Im[421], X_Im[420], X_Im[419], X_Im[418], X_Im[417], X_Im[416], X_Im[415], X_Im[414], X_Im[413], X_Im[412], X_Im[411], X_Im[410], X_Im[409], X_Im[408], X_Im[407], X_Im[406], X_Im[405], X_Im[404], X_Im[403], X_Im[402], X_Im[401], X_Im[400], X_Im[399], X_Im[398], X_Im[397], X_Im[396], X_Im[395], X_Im[394], X_Im[393], X_Im[392], X_Im[391], X_Im[390], X_Im[389], X_Im[388], X_Im[387], X_Im[386], X_Im[385], X_Im[384], X_Im[383], X_Im[382], X_Im[381], X_Im[380], X_Im[379], X_Im[378], X_Im[377], X_Im[376], X_Im[375], X_Im[374], X_Im[373], X_Im[372], X_Im[371], X_Im[370], X_Im[369], X_Im[368], X_Im[367], X_Im[366], X_Im[365], X_Im[364], X_Im[363], X_Im[362], X_Im[361], X_Im[360], X_Im[359], X_Im[358], X_Im[357], X_Im[356], X_Im[355], X_Im[354], X_Im[353], X_Im[352], X_Im[351], X_Im[350], X_Im[349], X_Im[348], X_Im[347], X_Im[346], X_Im[345], X_Im[344], X_Im[343], X_Im[342], X_Im[341], X_Im[340], X_Im[339], X_Im[338], X_Im[337], X_Im[336], X_Im[335], X_Im[334], X_Im[333], X_Im[332], X_Im[331], X_Im[330], X_Im[329], X_Im[328], X_Im[327], X_Im[326], X_Im[325], X_Im[324], X_Im[323], X_Im[322], X_Im[321], X_Im[320], X_Im[319], X_Im[318], X_Im[317], X_Im[316], X_Im[315], X_Im[314], X_Im[313], X_Im[312], X_Im[311], X_Im[310], X_Im[309], X_Im[308], X_Im[307], X_Im[306], X_Im[305], X_Im[304], X_Im[303], X_Im[302], X_Im[301], X_Im[300], X_Im[299], X_Im[298], X_Im[297], X_Im[296], X_Im[295], X_Im[294], X_Im[293], X_Im[292], X_Im[291], X_Im[290], X_Im[289], X_Im[288], X_Im[287], X_Im[286], X_Im[285], X_Im[284], X_Im[283], X_Im[282], X_Im[281], X_Im[280], X_Im[279], X_Im[278], X_Im[277], X_Im[276], X_Im[275], X_Im[274], X_Im[273], X_Im[272], X_Im[271], X_Im[270], X_Im[269], X_Im[268], X_Im[267], X_Im[266], X_Im[265], X_Im[264], X_Im[263], X_Im[262], X_Im[261], X_Im[260], X_Im[259], X_Im[258], X_Im[257], X_Im[256], X_Im[255], X_Im[254], X_Im[253], X_Im[252], X_Im[251], X_Im[250], X_Im[249], X_Im[248], X_Im[247], X_Im[246], X_Im[245], X_Im[244], X_Im[243], X_Im[242], X_Im[241], X_Im[240], X_Im[239], X_Im[238], X_Im[237], X_Im[236], X_Im[235], X_Im[234], X_Im[233], X_Im[232], X_Im[231], X_Im[230], X_Im[229], X_Im[228], X_Im[227], X_Im[226], X_Im[225], X_Im[224], X_Im[223], X_Im[222], X_Im[221], X_Im[220], X_Im[219], X_Im[218], X_Im[217], X_Im[216], X_Im[215], X_Im[214], X_Im[213], X_Im[212], X_Im[211], X_Im[210], X_Im[209], X_Im[208], X_Im[207], X_Im[206], X_Im[205], X_Im[204], X_Im[203], X_Im[202], X_Im[201], X_Im[200], X_Im[199], X_Im[198], X_Im[197], X_Im[196], X_Im[195], X_Im[194], X_Im[193], X_Im[192], X_Im[191], X_Im[190], X_Im[189], X_Im[188], X_Im[187], X_Im[186], X_Im[185], X_Im[184], X_Im[183], X_Im[182], X_Im[181], X_Im[180], X_Im[179], X_Im[178], X_Im[177], X_Im[176], X_Im[175], X_Im[174], X_Im[173], X_Im[172], X_Im[171], X_Im[170], X_Im[169], X_Im[168], X_Im[167], X_Im[166], X_Im[165], X_Im[164], X_Im[163], X_Im[162], X_Im[161], X_Im[160], X_Im[159], X_Im[158], X_Im[157], X_Im[156], X_Im[155], X_Im[154], X_Im[153], X_Im[152], X_Im[151], X_Im[150], X_Im[149], X_Im[148], X_Im[147], X_Im[146], X_Im[145], X_Im[144], X_Im[143], X_Im[142], X_Im[141], X_Im[140], X_Im[139], X_Im[138], X_Im[137], X_Im[136], X_Im[135], X_Im[134], X_Im[133], X_Im[132], X_Im[131], X_Im[130], X_Im[129], X_Im[128], X_Im[127], X_Im[126], X_Im[125], X_Im[124], X_Im[123], X_Im[122], X_Im[121], X_Im[120], X_Im[119], X_Im[118], X_Im[117], X_Im[116], X_Im[115], X_Im[114], X_Im[113], X_Im[112], X_Im[111], X_Im[110], X_Im[109], X_Im[108], X_Im[107], X_Im[106], X_Im[105], X_Im[104], X_Im[103], X_Im[102], X_Im[101], X_Im[100], X_Im[99], X_Im[98], X_Im[97], X_Im[96], X_Im[95], X_Im[94], X_Im[93], X_Im[92], X_Im[91], X_Im[90], X_Im[89], X_Im[88], X_Im[87], X_Im[86], X_Im[85], X_Im[84], X_Im[83], X_Im[82], X_Im[81], X_Im[80], X_Im[79], X_Im[78], X_Im[77], X_Im[76], X_Im[75], X_Im[74], X_Im[73], X_Im[72], X_Im[71], X_Im[70], X_Im[69], X_Im[68], X_Im[67], X_Im[66], X_Im[65], X_Im[64], X_Im[63], X_Im[62], X_Im[61], X_Im[60], X_Im[59], X_Im[58], X_Im[57], X_Im[56], X_Im[55], X_Im[54], X_Im[53], X_Im[52], X_Im[51], X_Im[50], X_Im[49], X_Im[48], X_Im[47], X_Im[46], X_Im[45], X_Im[44], X_Im[43], X_Im[42], X_Im[41], X_Im[40], X_Im[39], X_Im[38], X_Im[37], X_Im[36], X_Im[35], X_Im[34], X_Im[33], X_Im[32], X_Im[31], X_Im[30], X_Im[29], X_Im[28], X_Im[27], X_Im[26], X_Im[25], X_Im[24], X_Im[23], X_Im[22], X_Im[21], X_Im[20], X_Im[19], X_Im[18], X_Im[17], X_Im[16], X_Im[15], X_Im[14], X_Im[13], X_Im[12], X_Im[11], X_Im[10], X_Im[9], X_Im[8], X_Im[7], X_Im[6], X_Im[5], X_Im[4], X_Im[3], X_Im[2], X_Im[1], X_Im[0]};
	
	// Instantiate the Unit Under Test (UUT)
	FFT1024 uut (
		.Clk(Clk),
		.Reset(Reset),
		.Start(Start),
		.Ack(Ack),
		.x_re_packed(X_Re_Packed),
		.x_im_packed(32768'd0),
		.Done(Done),
		.state(state),
		.y_re_packed(Y_Re_out),
		.y_im_packed(Y_Im_out)
	);
	
	
	initial
	begin
		Clk = 0; // Initialize clock
		Start = 0;
		Reset = 0;
	end
	
	// Keep clock running
	always
	begin
		#20; 
		Clk = ~ Clk; 
	end
	
	initial
	begin
		Start = 0;
		Reset = 0;
		Ack = 0;
		#10
		Reset = 1;
		#200
		// FFT
X_Re[0]=32'd0; X_Re[1]=-32'd202; X_Re[2]=-32'd2459; X_Re[3]=-32'd1021; X_Re[4]=32'd202; X_Re[5]=32'd1248; X_Re[6]=32'd618; X_Re[7]=-32'd820; X_Re[8]=-32'd1021; X_Re[9]=-32'd2459; X_Re[10]=-32'd4123; X_Re[11]=-32'd4728; X_Re[12]=-32'd5939; X_Re[13]=-32'd6241; X_Re[14]=-32'd2459; X_Re[15]=-32'd416; X_Re[16]=-32'd1248; X_Re[17]=-32'd2459; X_Re[18]=32'd0; X_Re[19]=32'd2459; X_Re[20]=32'd4123; X_Re[21]=32'd5939; X_Re[22]=32'd4930; X_Re[23]=32'd4123; X_Re[24]=32'd2660; X_Re[25]=32'd1853; X_Re[26]=32'd0; X_Re[27]=-32'd2055; X_Re[28]=-32'd3114; X_Re[29]=-32'd1248; X_Re[30]=-32'd202; X_Re[31]=-32'd618; X_Re[32]=-32'd2459; X_Re[33]=-32'd3114; X_Re[34]=-32'd2459; X_Re[35]=-32'd2459; X_Re[36]=-32'd1021; X_Re[37]=-32'd1853; X_Re[38]=-32'd618; X_Re[39]=32'd820; X_Re[40]=32'd1853; X_Re[41]=32'd1853; X_Re[42]=32'd820; X_Re[43]=-32'd618; X_Re[44]=32'd820; X_Re[45]=32'd3518; X_Re[46]=32'd4123; X_Re[47]=32'd2660; X_Re[48]=32'd1021; X_Re[49]=32'd202; X_Re[50]=-32'd1021; X_Re[51]=32'd202; X_Re[52]=-32'd202; X_Re[53]=32'd820; X_Re[54]=32'd3921; X_Re[55]=32'd4930; X_Re[56]=32'd5334; X_Re[57]=32'd5334; X_Re[58]=32'd1652; X_Re[59]=32'd0; X_Re[60]=32'd202; X_Re[61]=-32'd202; X_Re[62]=-32'd3114; X_Re[63]=-32'd4123; X_Re[64]=-32'd4123; X_Re[65]=-32'd3720; X_Re[66]=-32'd1652; X_Re[67]=-32'd202; X_Re[68]=-32'd618; X_Re[69]=32'd618; X_Re[70]=32'd2660; X_Re[71]=32'd4728; X_Re[72]=32'd4930; X_Re[73]=32'd3518; X_Re[74]=32'd1652; X_Re[75]=32'd1853; X_Re[76]=32'd3921; X_Re[77]=32'd2459; X_Re[78]=32'd820; X_Re[79]=-32'd416; X_Re[80]=32'd618; X_Re[81]=32'd820; X_Re[82]=32'd1853; X_Re[83]=32'd1853; X_Re[84]=32'd1652; X_Re[85]=32'd820; X_Re[86]=-32'd202; X_Re[87]=-32'd820; X_Re[88]=-32'd1652; X_Re[89]=-32'd4728; X_Re[90]=-32'd3316; X_Re[91]=32'd1450; X_Re[92]=32'd2257; X_Re[93]=32'd1021; X_Re[94]=-32'd202; X_Re[95]=32'd0; X_Re[96]=32'd0; X_Re[97]=32'd2055; X_Re[98]=32'd3114; X_Re[99]=32'd2660; X_Re[100]=32'd3114; X_Re[101]=32'd2257; X_Re[102]=32'd1248; X_Re[103]=32'd618; X_Re[104]=-32'd3114; X_Re[105]=-32'd3518; X_Re[106]=-32'd618; X_Re[107]=32'd1652; X_Re[108]=32'd1652; X_Re[109]=32'd1450; X_Re[110]=32'd416; X_Re[111]=-32'd1853; X_Re[112]=-32'd2257; X_Re[113]=-32'd2459; X_Re[114]=-32'd2660; X_Re[115]=-32'd2459; X_Re[116]=-32'd3518; X_Re[117]=-32'd2913; X_Re[118]=-32'd2257; X_Re[119]=-32'd3316; X_Re[120]=-32'd4930; X_Re[121]=-32'd2459; X_Re[122]=32'd1853; X_Re[123]=32'd2913; X_Re[124]=32'd4123; X_Re[125]=32'd3921; X_Re[126]=32'd1853; X_Re[127]=32'd820; X_Re[128]=32'd2257; X_Re[129]=32'd1652; X_Re[130]=32'd820; X_Re[131]=32'd618; X_Re[132]=32'd1021; X_Re[133]=32'd1652; X_Re[134]=32'd416; X_Re[135]=-32'd2055; X_Re[136]=-32'd2660; X_Re[137]=-32'd2660; X_Re[138]=-32'd3518; X_Re[139]=-32'd3114; X_Re[140]=-32'd3518; X_Re[141]=-32'd3518; X_Re[142]=-32'd3114; X_Re[143]=-32'd202; X_Re[144]=32'd202; X_Re[145]=32'd416; X_Re[146]=32'd1853; X_Re[147]=32'd1853; X_Re[148]=32'd1853; X_Re[149]=32'd2257; X_Re[150]=32'd820; X_Re[151]=-32'd820; X_Re[152]=32'd618; X_Re[153]=32'd1248; X_Re[154]=32'd820; X_Re[155]=-32'd202; X_Re[156]=-32'd618; X_Re[157]=-32'd618; X_Re[158]=32'd1021; X_Re[159]=32'd3114; X_Re[160]=32'd3114; X_Re[161]=32'd3720; X_Re[162]=32'd1248; X_Re[163]=-32'd416; X_Re[164]=-32'd1652; X_Re[165]=-32'd5132; X_Re[166]=-32'd7452; X_Re[167]=-32'd6241; X_Re[168]=-32'd3720; X_Re[169]=-32'd2257; X_Re[170]=-32'd202; X_Re[171]=32'd202; X_Re[172]=-32'd416; X_Re[173]=32'd1450; X_Re[174]=32'd3921; X_Re[175]=32'd4325; X_Re[176]=32'd4930; X_Re[177]=32'd5132; X_Re[178]=32'd4123; X_Re[179]=32'd3518; X_Re[180]=32'd1248; X_Re[181]=-32'd1652; X_Re[182]=-32'd3518; X_Re[183]=-32'd1652; X_Re[184]=32'd618; X_Re[185]=32'd1021; X_Re[186]=32'd1652; X_Re[187]=32'd0; X_Re[188]=-32'd1248; X_Re[189]=-32'd1450; X_Re[190]=-32'd2055; X_Re[191]=-32'd1450; X_Re[192]=-32'd202; X_Re[193]=32'd0; X_Re[194]=32'd416; X_Re[195]=32'd820; X_Re[196]=-32'd618; X_Re[197]=-32'd1652; X_Re[198]=-32'd618; X_Re[199]=32'd1021; X_Re[200]=32'd1652; X_Re[201]=32'd3720; X_Re[202]=32'd2913; X_Re[203]=32'd1248; X_Re[204]=32'd1021; X_Re[205]=32'd1450; X_Re[206]=32'd1021; X_Re[207]=32'd820; X_Re[208]=32'd1450; X_Re[209]=32'd1853; X_Re[210]=32'd2660; X_Re[211]=32'd2055; X_Re[212]=32'd1021; X_Re[213]=-32'd202; X_Re[214]=-32'd416; X_Re[215]=-32'd618; X_Re[216]=-32'd416; X_Re[217]=-32'd1853; X_Re[218]=-32'd3921; X_Re[219]=-32'd4123; X_Re[220]=-32'd3921; X_Re[221]=-32'd3921; X_Re[222]=-32'd2459; X_Re[223]=-32'd1021; X_Re[224]=-32'd1450; X_Re[225]=-32'd416; X_Re[226]=32'd618; X_Re[227]=32'd618; X_Re[228]=32'd1021; X_Re[229]=32'd2660; X_Re[230]=32'd4527; X_Re[231]=32'd4728; X_Re[232]=32'd4123; X_Re[233]=32'd416; X_Re[234]=-32'd820; X_Re[235]=-32'd416; X_Re[236]=32'd416; X_Re[237]=32'd202; X_Re[238]=32'd1021; X_Re[239]=32'd202; X_Re[240]=-32'd1853; X_Re[241]=-32'd4325; X_Re[242]=-32'd5334; X_Re[243]=-32'd5535; X_Re[244]=-32'd4728; X_Re[245]=-32'd2660; X_Re[246]=-32'd202; X_Re[247]=32'd1450; X_Re[248]=32'd1450; X_Re[249]=32'd1021; X_Re[250]=32'd1652; X_Re[251]=32'd1248; X_Re[252]=32'd1021; X_Re[253]=32'd2257; X_Re[254]=32'd2660; X_Re[255]=32'd820; X_Re[256]=32'd0; X_Re[257]=-32'd1021; X_Re[258]=-32'd3114; X_Re[259]=-32'd3316; X_Re[260]=32'd416; X_Re[261]=32'd2459; X_Re[262]=32'd4123; X_Re[263]=32'd3921; X_Re[264]=32'd2459; X_Re[265]=32'd1248; X_Re[266]=32'd0; X_Re[267]=-32'd1652; X_Re[268]=-32'd2257; X_Re[269]=-32'd2257; X_Re[270]=-32'd3114; X_Re[271]=-32'd3720; X_Re[272]=-32'd3518; X_Re[273]=-32'd3921; X_Re[274]=-32'd3720; X_Re[275]=-32'd1450; X_Re[276]=32'd1021; X_Re[277]=32'd3720; X_Re[278]=32'd4728; X_Re[279]=32'd3720; X_Re[280]=32'd3316; X_Re[281]=32'd4123; X_Re[282]=32'd3316; X_Re[283]=32'd3114; X_Re[284]=32'd2913; X_Re[285]=32'd1248; X_Re[286]=32'd618; X_Re[287]=32'd820; X_Re[288]=32'd820; X_Re[289]=-32'd618; X_Re[290]=-32'd1021; X_Re[291]=-32'd618; X_Re[292]=-32'd416; X_Re[293]=32'd202; X_Re[294]=-32'd416; X_Re[295]=-32'd1450; X_Re[296]=-32'd2055; X_Re[297]=-32'd1853; X_Re[298]=-32'd1248; X_Re[299]=32'd618; X_Re[300]=32'd820; X_Re[301]=32'd820; X_Re[302]=-32'd416; X_Re[303]=-32'd202; X_Re[304]=-32'd820; X_Re[305]=-32'd202; X_Re[306]=32'd1652; X_Re[307]=32'd3114; X_Re[308]=32'd3921; X_Re[309]=32'd2660; X_Re[310]=32'd202; X_Re[311]=-32'd416; X_Re[312]=32'd1021; X_Re[313]=32'd1021; X_Re[314]=32'd1021; X_Re[315]=32'd3114; X_Re[316]=32'd2257; X_Re[317]=-32'd202; X_Re[318]=-32'd1248; X_Re[319]=-32'd2660; X_Re[320]=-32'd4728; X_Re[321]=-32'd4325; X_Re[322]=-32'd2660; X_Re[323]=-32'd1450; X_Re[324]=-32'd1652; X_Re[325]=-32'd1248; X_Re[326]=-32'd1021; X_Re[327]=-32'd202; X_Re[328]=-32'd820; X_Re[329]=32'd416; X_Re[330]=32'd1652; X_Re[331]=32'd1853; X_Re[332]=32'd2055; X_Re[333]=32'd1853; X_Re[334]=32'd0; X_Re[335]=-32'd2660; X_Re[336]=-32'd2913; X_Re[337]=-32'd1021; X_Re[338]=32'd1248; X_Re[339]=32'd1450; X_Re[340]=32'd820; X_Re[341]=32'd202; X_Re[342]=-32'd1021; X_Re[343]=-32'd2913; X_Re[344]=-32'd2660; X_Re[345]=-32'd1853; X_Re[346]=-32'd1450; X_Re[347]=-32'd2257; X_Re[348]=-32'd2660; X_Re[349]=-32'd3114; X_Re[350]=-32'd3518; X_Re[351]=-32'd2660; X_Re[352]=32'd0; X_Re[353]=32'd1652; X_Re[354]=32'd2257; X_Re[355]=32'd1652; X_Re[356]=32'd1021; X_Re[357]=32'd1450; X_Re[358]=32'd1450; X_Re[359]=32'd1021; X_Re[360]=32'd618; X_Re[361]=32'd618; X_Re[362]=32'd416; X_Re[363]=32'd1021; X_Re[364]=32'd2055; X_Re[365]=32'd1021; X_Re[366]=32'd618; X_Re[367]=32'd2257; X_Re[368]=32'd3114; X_Re[369]=32'd3518; X_Re[370]=32'd1853; X_Re[371]=-32'd202; X_Re[372]=-32'd1853; X_Re[373]=-32'd3316; X_Re[374]=-32'd4728; X_Re[375]=-32'd4123; X_Re[376]=-32'd2913; X_Re[377]=-32'd1853; X_Re[378]=-32'd2257; X_Re[379]=-32'd2257; X_Re[380]=-32'd1450; X_Re[381]=-32'd1248; X_Re[382]=32'd820; X_Re[383]=32'd4527; X_Re[384]=32'd7452; X_Re[385]=32'd7048; X_Re[386]=32'd5132; X_Re[387]=32'd3316; X_Re[388]=32'd1853; X_Re[389]=32'd1021; X_Re[390]=32'd820; X_Re[391]=32'd1450; X_Re[392]=32'd1248; X_Re[393]=-32'd1450; X_Re[394]=-32'd2257; X_Re[395]=-32'd2660; X_Re[396]=-32'd4325; X_Re[397]=-32'd3921; X_Re[398]=-32'd1853; X_Re[399]=32'd618; X_Re[400]=32'd0; X_Re[401]=32'd820; X_Re[402]=32'd2055; X_Re[403]=32'd2055; X_Re[404]=32'd1450; X_Re[405]=32'd1248; X_Re[406]=32'd1450; X_Re[407]=32'd1652; X_Re[408]=32'd618; X_Re[409]=32'd1248; X_Re[410]=32'd820; X_Re[411]=-32'd1652; X_Re[412]=-32'd2257; X_Re[413]=32'd202; X_Re[414]=32'd3114; X_Re[415]=32'd3921; X_Re[416]=32'd3720; X_Re[417]=32'd3518; X_Re[418]=32'd2257; X_Re[419]=32'd820; X_Re[420]=-32'd416; X_Re[421]=-32'd618; X_Re[422]=-32'd820; X_Re[423]=-32'd2055; X_Re[424]=-32'd2660; X_Re[425]=-32'd3316; X_Re[426]=-32'd4930; X_Re[427]=-32'd4930; X_Re[428]=-32'd2459; X_Re[429]=-32'd618; X_Re[430]=32'd1248; X_Re[431]=32'd820; X_Re[432]=32'd2459; X_Re[433]=32'd3114; X_Re[434]=32'd2913; X_Re[435]=32'd2459; X_Re[436]=32'd2459; X_Re[437]=32'd1450; X_Re[438]=32'd1021; X_Re[439]=32'd0; X_Re[440]=-32'd202; X_Re[441]=-32'd618; X_Re[442]=-32'd416; X_Re[443]=32'd416; X_Re[444]=32'd1652; X_Re[445]=32'd2660; X_Re[446]=32'd1450; X_Re[447]=32'd618; X_Re[448]=32'd0; X_Re[449]=-32'd416; X_Re[450]=-32'd1652; X_Re[451]=-32'd3720; X_Re[452]=-32'd3921; X_Re[453]=-32'd2913; X_Re[454]=-32'd3114; X_Re[455]=-32'd2459; X_Re[456]=-32'd2055; X_Re[457]=-32'd2913; X_Re[458]=-32'd2257; X_Re[459]=32'd1021; X_Re[460]=32'd4325; X_Re[461]=32'd4527; X_Re[462]=32'd2913; X_Re[463]=32'd2055; X_Re[464]=32'd1652; X_Re[465]=32'd618; X_Re[466]=-32'd202; X_Re[467]=32'd1450; X_Re[468]=32'd1853; X_Re[469]=32'd416; X_Re[470]=-32'd820; X_Re[471]=-32'd202; X_Re[472]=-32'd2055; X_Re[473]=-32'd3114; X_Re[474]=-32'd2055; X_Re[475]=-32'd416; X_Re[476]=-32'd618; X_Re[477]=-32'd1652; X_Re[478]=-32'd1248; X_Re[479]=-32'd1450; X_Re[480]=-32'd2257; X_Re[481]=-32'd2660; X_Re[482]=-32'd1853; X_Re[483]=-32'd1450; X_Re[484]=-32'd1021; X_Re[485]=-32'd416; X_Re[486]=32'd820; X_Re[487]=32'd416; X_Re[488]=-32'd820; X_Re[489]=32'd618; X_Re[490]=32'd2660; X_Re[491]=32'd3316; X_Re[492]=32'd2913; X_Re[493]=32'd2913; X_Re[494]=32'd2055; X_Re[495]=32'd416; X_Re[496]=-32'd1021; X_Re[497]=-32'd1853; X_Re[498]=-32'd1853; X_Re[499]=-32'd1853; X_Re[500]=-32'd2055; X_Re[501]=-32'd1450; X_Re[502]=-32'd1853; X_Re[503]=-32'd3114; X_Re[504]=-32'd1853; X_Re[505]=-32'd202; X_Re[506]=32'd1450; X_Re[507]=32'd1450; X_Re[508]=32'd416; X_Re[509]=32'd416; X_Re[510]=32'd416; X_Re[511]=32'd618; X_Re[512]=32'd202; X_Re[513]=-32'd202; X_Re[514]=-32'd202; X_Re[515]=32'd0; X_Re[516]=-32'd202; X_Re[517]=32'd416; X_Re[518]=32'd618; X_Re[519]=32'd1853; X_Re[520]=32'd3921; X_Re[521]=32'd5334; X_Re[522]=32'd4527; X_Re[523]=32'd3720; X_Re[524]=32'd2660; X_Re[525]=32'd1450; X_Re[526]=-32'd618; X_Re[527]=-32'd2257; X_Re[528]=-32'd4123; X_Re[529]=-32'd4123; X_Re[530]=-32'd4527; X_Re[531]=-32'd4527; X_Re[532]=-32'd3720; X_Re[533]=-32'd2459; X_Re[534]=-32'd1652; X_Re[535]=32'd1652; X_Re[536]=32'd3921; X_Re[537]=32'd6241; X_Re[538]=32'd5535; X_Re[539]=32'd4728; X_Re[540]=32'd4527; X_Re[541]=32'd3921; X_Re[542]=32'd2257; X_Re[543]=32'd1021; X_Re[544]=32'd820; X_Re[545]=32'd0; X_Re[546]=-32'd820; X_Re[547]=-32'd820; X_Re[548]=-32'd1450; X_Re[549]=-32'd2055; X_Re[550]=-32'd1248; X_Re[551]=32'd1248; X_Re[552]=32'd2660; X_Re[553]=32'd1450; X_Re[554]=32'd1248; X_Re[555]=32'd820; X_Re[556]=32'd618; X_Re[557]=32'd0; X_Re[558]=-32'd202; X_Re[559]=-32'd618; X_Re[560]=-32'd1021; X_Re[561]=-32'd1248; X_Re[562]=-32'd618; X_Re[563]=-32'd202; X_Re[564]=-32'd416; X_Re[565]=-32'd618; X_Re[566]=32'd1021; X_Re[567]=32'd1853; X_Re[568]=32'd2055; X_Re[569]=32'd2257; X_Re[570]=32'd2257; X_Re[571]=32'd2055; X_Re[572]=32'd1248; X_Re[573]=-32'd202; X_Re[574]=-32'd1450; X_Re[575]=-32'd1652; X_Re[576]=-32'd2055; X_Re[577]=-32'd2660; X_Re[578]=-32'd2913; X_Re[579]=-32'd3114; X_Re[580]=-32'd3316; X_Re[581]=-32'd2660; X_Re[582]=-32'd618; X_Re[583]=-32'd416; X_Re[584]=-32'd618; X_Re[585]=32'd0; X_Re[586]=32'd820; X_Re[587]=32'd1450; X_Re[588]=32'd1450; X_Re[589]=32'd1248; X_Re[590]=32'd0; X_Re[591]=32'd0; X_Re[592]=-32'd618; X_Re[593]=-32'd820; X_Re[594]=-32'd820; X_Re[595]=-32'd1021; X_Re[596]=32'd202; X_Re[597]=32'd1652; X_Re[598]=32'd2257; X_Re[599]=32'd1450; X_Re[600]=32'd618; X_Re[601]=32'd1021; X_Re[602]=32'd1021; X_Re[603]=32'd202; X_Re[604]=-32'd1021; X_Re[605]=-32'd2257; X_Re[606]=-32'd2913; X_Re[607]=-32'd3316; X_Re[608]=-32'd2459; X_Re[609]=-32'd2660; X_Re[610]=-32'd2459; X_Re[611]=-32'd1652; X_Re[612]=-32'd416; X_Re[613]=32'd1450; X_Re[614]=32'd2055; X_Re[615]=32'd1853; X_Re[616]=32'd2257; X_Re[617]=32'd2660; X_Re[618]=32'd1853; X_Re[619]=32'd820; X_Re[620]=32'd202; X_Re[621]=32'd0; X_Re[622]=-32'd202; X_Re[623]=-32'd202; X_Re[624]=32'd0; X_Re[625]=-32'd618; X_Re[626]=-32'd618; X_Re[627]=32'd820; X_Re[628]=32'd1652; X_Re[629]=32'd1450; X_Re[630]=32'd618; X_Re[631]=-32'd618; X_Re[632]=-32'd1021; X_Re[633]=-32'd1248; X_Re[634]=-32'd1450; X_Re[635]=-32'd2913; X_Re[636]=-32'd3720; X_Re[637]=-32'd2913; X_Re[638]=-32'd1853; X_Re[639]=-32'd618; X_Re[640]=32'd820; X_Re[641]=32'd1021; X_Re[642]=32'd2257; X_Re[643]=32'd3114; X_Re[644]=32'd3114; X_Re[645]=32'd2459; X_Re[646]=32'd2055; X_Re[647]=32'd1853; X_Re[648]=32'd1450; X_Re[649]=32'd1021; X_Re[650]=32'd0; X_Re[651]=-32'd1652; X_Re[652]=-32'd2055; X_Re[653]=-32'd1450; X_Re[654]=-32'd1021; X_Re[655]=-32'd1021; X_Re[656]=-32'd618; X_Re[657]=-32'd416; X_Re[658]=-32'd416; X_Re[659]=32'd618; X_Re[660]=32'd1248; X_Re[661]=32'd820; X_Re[662]=32'd1450; X_Re[663]=32'd1021; X_Re[664]=32'd618; X_Re[665]=32'd202; X_Re[666]=-32'd202; X_Re[667]=-32'd1021; X_Re[668]=-32'd416; X_Re[669]=-32'd202; X_Re[670]=-32'd416; X_Re[671]=32'd618; X_Re[672]=32'd2257; X_Re[673]=32'd3720; X_Re[674]=32'd4527; X_Re[675]=32'd5132; X_Re[676]=32'd4325; X_Re[677]=32'd3921; X_Re[678]=32'd3720; X_Re[679]=32'd2660; X_Re[680]=32'd202; X_Re[681]=-32'd2055; X_Re[682]=-32'd4325; X_Re[683]=-32'd5132; X_Re[684]=-32'd5535; X_Re[685]=-32'd4930; X_Re[686]=-32'd4325; X_Re[687]=-32'd3720; X_Re[688]=-32'd2055; X_Re[689]=-32'd416; X_Re[690]=32'd1021; X_Re[691]=32'd1853; X_Re[692]=32'd2459; X_Re[693]=32'd3720; X_Re[694]=32'd4728; X_Re[695]=32'd3518; X_Re[696]=32'd2257; X_Re[697]=-32'd202; X_Re[698]=-32'd1248; X_Re[699]=-32'd2257; X_Re[700]=-32'd2257; X_Re[701]=-32'd2660; X_Re[702]=-32'd2257; X_Re[703]=-32'd1652; X_Re[704]=-32'd202; X_Re[705]=32'd618; X_Re[706]=32'd820; X_Re[707]=32'd618; X_Re[708]=32'd1248; X_Re[709]=32'd1248; X_Re[710]=32'd202; X_Re[711]=-32'd618; X_Re[712]=-32'd2459; X_Re[713]=-32'd3316; X_Re[714]=-32'd3316; X_Re[715]=-32'd3114; X_Re[716]=-32'd2913; X_Re[717]=-32'd1652; X_Re[718]=-32'd618; X_Re[719]=32'd820; X_Re[720]=32'd2055; X_Re[721]=32'd2459; X_Re[722]=32'd2055; X_Re[723]=32'd2055; X_Re[724]=32'd2660; X_Re[725]=32'd2913; X_Re[726]=32'd2257; X_Re[727]=32'd1021; X_Re[728]=-32'd618; X_Re[729]=-32'd820; X_Re[730]=-32'd820; X_Re[731]=-32'd1021; X_Re[732]=-32'd820; X_Re[733]=-32'd416; X_Re[734]=-32'd1021; X_Re[735]=-32'd1248; X_Re[736]=-32'd1248; X_Re[737]=-32'd618; X_Re[738]=-32'd416; X_Re[739]=32'd202; X_Re[740]=32'd1021; X_Re[741]=32'd1021; X_Re[742]=-32'd202; X_Re[743]=-32'd820; X_Re[744]=32'd0; X_Re[745]=32'd202; X_Re[746]=32'd820; X_Re[747]=32'd820; X_Re[748]=32'd1450; X_Re[749]=32'd1021; X_Re[750]=32'd1450; X_Re[751]=32'd2055; X_Re[752]=32'd2257; X_Re[753]=32'd2913; X_Re[754]=32'd3316; X_Re[755]=32'd3518; X_Re[756]=32'd2459; X_Re[757]=32'd618; X_Re[758]=-32'd820; X_Re[759]=-32'd2459; X_Re[760]=-32'd3114; X_Re[761]=-32'd3316; X_Re[762]=-32'd2913; X_Re[763]=-32'd1853; X_Re[764]=-32'd416; X_Re[765]=32'd202; X_Re[766]=32'd416; X_Re[767]=32'd618; X_Re[768]=32'd618; X_Re[769]=32'd1853; X_Re[770]=32'd3316; X_Re[771]=32'd3518; X_Re[772]=32'd2913; X_Re[773]=32'd618; X_Re[774]=-32'd1248; X_Re[775]=-32'd1450; X_Re[776]=-32'd820; X_Re[777]=-32'd820; X_Re[778]=-32'd416; X_Re[779]=32'd1021; X_Re[780]=32'd1450; X_Re[781]=32'd1853; X_Re[782]=32'd2055; X_Re[783]=32'd1652; X_Re[784]=32'd1450; X_Re[785]=32'd1248; X_Re[786]=32'd202; X_Re[787]=-32'd1021; X_Re[788]=-32'd2459; X_Re[789]=-32'd3316; X_Re[790]=-32'd3518; X_Re[791]=-32'd2913; X_Re[792]=-32'd2459; X_Re[793]=-32'd2055; X_Re[794]=-32'd1450; X_Re[795]=32'd0; X_Re[796]=32'd1021; X_Re[797]=32'd2055; X_Re[798]=32'd2660; X_Re[799]=32'd2257; X_Re[800]=32'd1450; X_Re[801]=32'd1652; X_Re[802]=32'd1021; X_Re[803]=-32'd820; X_Re[804]=-32'd2660; X_Re[805]=-32'd2660; X_Re[806]=-32'd3114; X_Re[807]=-32'd2257; X_Re[808]=-32'd1652; X_Re[809]=-32'd1021; X_Re[810]=32'd202; X_Re[811]=32'd416; X_Re[812]=-32'd202; X_Re[813]=32'd202; X_Re[814]=32'd416; X_Re[815]=32'd416; X_Re[816]=32'd820; X_Re[817]=32'd618; X_Re[818]=-32'd1021; X_Re[819]=-32'd3114; X_Re[820]=-32'd3518; X_Re[821]=-32'd3518; X_Re[822]=-32'd1853; X_Re[823]=-32'd618; X_Re[824]=32'd618; X_Re[825]=32'd1021; X_Re[826]=32'd1450; X_Re[827]=32'd1853; X_Re[828]=32'd2055; X_Re[829]=32'd2055; X_Re[830]=32'd2459; X_Re[831]=32'd3316; X_Re[832]=32'd3316; X_Re[833]=32'd2459; X_Re[834]=32'd1021; X_Re[835]=-32'd1021; X_Re[836]=-32'd2055; X_Re[837]=-32'd2660; X_Re[838]=-32'd3518; X_Re[839]=-32'd3316; X_Re[840]=-32'd1652; X_Re[841]=-32'd202; X_Re[842]=32'd202; X_Re[843]=32'd416; X_Re[844]=32'd1021; X_Re[845]=32'd1652; X_Re[846]=32'd2660; X_Re[847]=32'd3316; X_Re[848]=32'd4527; X_Re[849]=32'd3316; X_Re[850]=32'd1450; X_Re[851]=-32'd202; X_Re[852]=-32'd1652; X_Re[853]=-32'd1450; X_Re[854]=-32'd1853; X_Re[855]=-32'd1248; X_Re[856]=32'd0; X_Re[857]=32'd1021; X_Re[858]=32'd1248; X_Re[859]=32'd2660; X_Re[860]=32'd2660; X_Re[861]=32'd2660; X_Re[862]=32'd3518; X_Re[863]=32'd2257; X_Re[864]=-32'd202; X_Re[865]=-32'd1652; X_Re[866]=-32'd2055; X_Re[867]=-32'd2257; X_Re[868]=-32'd1652; X_Re[869]=-32'd1652; X_Re[870]=-32'd1450; X_Re[871]=-32'd1021; X_Re[872]=-32'd820; X_Re[873]=-32'd820; X_Re[874]=32'd202; X_Re[875]=32'd1450; X_Re[876]=32'd1248; X_Re[877]=32'd1853; X_Re[878]=32'd2459; X_Re[879]=32'd1853; X_Re[880]=-32'd202; X_Re[881]=-32'd202; X_Re[882]=-32'd820; X_Re[883]=-32'd618; X_Re[884]=32'd416; X_Re[885]=32'd1021; X_Re[886]=32'd416; X_Re[887]=32'd820; X_Re[888]=32'd416; X_Re[889]=-32'd618; X_Re[890]=-32'd416; X_Re[891]=-32'd202; X_Re[892]=32'd416; X_Re[893]=32'd820; X_Re[894]=32'd618; X_Re[895]=-32'd1652; X_Re[896]=-32'd2459; X_Re[897]=-32'd3114; X_Re[898]=-32'd3114; X_Re[899]=-32'd1248; X_Re[900]=32'd1021; X_Re[901]=32'd1248; X_Re[902]=32'd2257; X_Re[903]=32'd2913; X_Re[904]=32'd2055; X_Re[905]=32'd2257; X_Re[906]=32'd2660; X_Re[907]=32'd2257; X_Re[908]=32'd2660; X_Re[909]=32'd3114; X_Re[910]=32'd1652; X_Re[911]=-32'd416; X_Re[912]=-32'd1450; X_Re[913]=-32'd2055; X_Re[914]=-32'd2913; X_Re[915]=-32'd2660; X_Re[916]=-32'd2913; X_Re[917]=-32'd2055; X_Re[918]=-32'd1450; X_Re[919]=-32'd1248; X_Re[920]=-32'd1021; X_Re[921]=-32'd416; X_Re[922]=-32'd202; X_Re[923]=32'd0; X_Re[924]=32'd820; X_Re[925]=32'd820; X_Re[926]=32'd202; X_Re[927]=32'd0; X_Re[928]=-32'd618; X_Re[929]=-32'd820; X_Re[930]=-32'd1248; X_Re[931]=-32'd1248; X_Re[932]=-32'd1021; X_Re[933]=-32'd202; X_Re[934]=32'd618; X_Re[935]=32'd1450; X_Re[936]=32'd2257; X_Re[937]=32'd2660; X_Re[938]=32'd2913; X_Re[939]=32'd2660; X_Re[940]=32'd1021; X_Re[941]=-32'd1021; X_Re[942]=-32'd3114; X_Re[943]=-32'd3720; X_Re[944]=-32'd3518; X_Re[945]=-32'd3518; X_Re[946]=-32'd2055; X_Re[947]=-32'd1853; X_Re[948]=-32'd202; X_Re[949]=32'd0; X_Re[950]=32'd0; X_Re[951]=32'd1248; X_Re[952]=32'd2257; X_Re[953]=32'd2660; X_Re[954]=32'd3720; X_Re[955]=32'd3720; X_Re[956]=32'd1450; X_Re[957]=-32'd618; X_Re[958]=-32'd1652; X_Re[959]=-32'd2459; X_Re[960]=-32'd1853; X_Re[961]=-32'd618; X_Re[962]=-32'd820; X_Re[963]=32'd618; X_Re[964]=32'd1652; X_Re[965]=32'd1021; X_Re[966]=32'd416; X_Re[967]=32'd618; X_Re[968]=32'd618; X_Re[969]=32'd820; X_Re[970]=32'd1652; X_Re[971]=32'd416; X_Re[972]=-32'd1021; X_Re[973]=-32'd2913; X_Re[974]=-32'd3114; X_Re[975]=-32'd3518; X_Re[976]=-32'd2913; X_Re[977]=-32'd1853; X_Re[978]=-32'd416; X_Re[979]=32'd1021; X_Re[980]=32'd1652; X_Re[981]=32'd1853; X_Re[982]=32'd2660; X_Re[983]=32'd2459; X_Re[984]=32'd2055; X_Re[985]=32'd2913; X_Re[986]=32'd2913; X_Re[987]=32'd618; X_Re[988]=-32'd1021; X_Re[989]=-32'd1248; X_Re[990]=-32'd1853; X_Re[991]=-32'd1853; X_Re[992]=-32'd1652; X_Re[993]=-32'd2257; X_Re[994]=-32'd1450; X_Re[995]=-32'd416; X_Re[996]=32'd0; X_Re[997]=32'd1248; X_Re[998]=32'd1853; X_Re[999]=32'd2055; X_Re[1000]=32'd2660; X_Re[1001]=32'd2055; X_Re[1002]=32'd820; X_Re[1003]=-32'd416; X_Re[1004]=-32'd1450; X_Re[1005]=-32'd1021; X_Re[1006]=-32'd1021; X_Re[1007]=-32'd618; X_Re[1008]=-32'd820; X_Re[1009]=-32'd618; X_Re[1010]=-32'd202; X_Re[1011]=32'd202; X_Re[1012]=32'd1021; X_Re[1013]=32'd1853; X_Re[1014]=32'd3114; X_Re[1015]=32'd3921; X_Re[1016]=32'd4123; X_Re[1017]=32'd2660; X_Re[1018]=32'd416; X_Re[1019]=-32'd1248; X_Re[1020]=-32'd1450; X_Re[1021]=-32'd1652; X_Re[1022]=-32'd1450; X_Re[1023]=-32'd1450;
		#10
		Reset = 0;
		#10
		
		Start = 1;
		//#32000
		#130
		Start = 0;
		Ack = 1;
		//$display("Results 1:");
		//$display("Y[0] expected %d+i%d got %d+i%d", -482739591, 0, Y_Re[0], Y_Im[0]);
		//$display("Y[1] expected %d+i%d got %d+i%d", 322112716, 107370905, Y_Re[1], Y_Im[1]);
		//$display("Y[2] expected %d+i%d got %d+i%d", -161485842, 0, Y_Re[2], Y_Im[2]);
		//$display("Y[3] expected %d+i%d got %d+i%d", 322112716, -107370905, Y_Re[3], Y_Im[3]);
		//#100
		//X_Re[0] = 16'd406;
		//X_Re[1] = 16'd2496;
		//X_Re[2] = 16'd1238;
		//X_Re[3] = -16'd1638;	  
		//#50
		//$display("Results 2:");
		//$display("Y[0] expected %d+i%d got %d+i%d", 164062743, 0, Y_Re[0], Y_Im[0]);
		//$display("Y[1] expected %d+i%d got %d+i%d", -054544420, 271004165, Y_Re[1], Y_Im[1]);
		//$display("Y[2] expected %d+i%d got %d+i%d", 051538034, 0, Y_Re[2], Y_Im[2]);
		//$display("Y[3] expected %d+i%d got %d+i%d", -054544420, -271004165, Y_Re[3], Y_Im[3]);
	end

endmodule