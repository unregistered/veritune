module FFT1024_LUT(n, twiddle);
	input [9:0] n;
		
	output reg [31:0] twiddle;
	
	always @ (n)
	begin
		//$display("LUT address=%d", n);
		case(n)
		8'd0  : twiddle = { 16'd32767   ,  16'd0       }; //i=0  n=256 twiddle= 1               + i 0
		8'd1  : twiddle = { 16'd32757   , -16'd804     }; //i=1  n=256 twiddle= 9.996988e-01    + i -2.454123e-02
		8'd2  : twiddle = { 16'd32728   , -16'd1608    }; //i=2  n=256 twiddle= 9.987955e-01    + i -4.906767e-02
		8'd3  : twiddle = { 16'd32678   , -16'd2410    }; //i=3  n=256 twiddle= 9.972905e-01    + i -7.356456e-02
		8'd4  : twiddle = { 16'd32609   , -16'd3212    }; //i=4  n=256 twiddle= 9.951847e-01    + i -9.801714e-02
		8'd5  : twiddle = { 16'd32521   , -16'd4011    }; //i=5  n=256 twiddle= 9.924795e-01    + i -1.224107e-01
		8'd6  : twiddle = { 16'd32412   , -16'd4808    }; //i=6  n=256 twiddle= 9.891765e-01    + i -1.467305e-01
		8'd7  : twiddle = { 16'd32285   , -16'd5602    }; //i=7  n=256 twiddle= 9.852776e-01    + i -1.709619e-01
		8'd8  : twiddle = { 16'd32137   , -16'd6393    }; //i=8  n=256 twiddle= 9.807853e-01    + i -1.950903e-01
		8'd9  : twiddle = { 16'd31971   , -16'd7179    }; //i=9  n=256 twiddle= 9.757021e-01    + i -2.191012e-01
		8'd10 : twiddle = { 16'd31785   , -16'd7962    }; //i=10 n=256 twiddle= 9.700313e-01    + i -2.429802e-01
		8'd11 : twiddle = { 16'd31580   , -16'd8739    }; //i=11 n=256 twiddle= 9.637761e-01    + i -2.667128e-01
		8'd12 : twiddle = { 16'd31356   , -16'd9512    }; //i=12 n=256 twiddle= 9.569403e-01    + i -2.902847e-01
		8'd13 : twiddle = { 16'd31113   , -16'd10278   }; //i=13 n=256 twiddle= 9.495282e-01    + i -3.136817e-01
		8'd14 : twiddle = { 16'd30852   , -16'd11039   }; //i=14 n=256 twiddle= 9.415441e-01    + i -3.368899e-01
		8'd15 : twiddle = { 16'd30571   , -16'd11793   }; //i=15 n=256 twiddle= 9.329928e-01    + i -3.598950e-01
		8'd16 : twiddle = { 16'd30273   , -16'd12539   }; //i=16 n=256 twiddle= 9.238795e-01    + i -3.826834e-01
		8'd17 : twiddle = { 16'd29956   , -16'd13279   }; //i=17 n=256 twiddle= 9.142098e-01    + i -4.052413e-01
		8'd18 : twiddle = { 16'd29621   , -16'd14010   }; //i=18 n=256 twiddle= 9.039893e-01    + i -4.275551e-01
		8'd19 : twiddle = { 16'd29268   , -16'd14732   }; //i=19 n=256 twiddle= 8.932243e-01    + i -4.496113e-01
		8'd20 : twiddle = { 16'd28898   , -16'd15446   }; //i=20 n=256 twiddle= 8.819213e-01    + i -4.713967e-01
		8'd21 : twiddle = { 16'd28510   , -16'd16151   }; //i=21 n=256 twiddle= 8.700870e-01    + i -4.928982e-01
		8'd22 : twiddle = { 16'd28105   , -16'd16846   }; //i=22 n=256 twiddle= 8.577286e-01    + i -5.141027e-01
		8'd23 : twiddle = { 16'd27683   , -16'd17530   }; //i=23 n=256 twiddle= 8.448536e-01    + i -5.349976e-01
		8'd24 : twiddle = { 16'd27245   , -16'd18204   }; //i=24 n=256 twiddle= 8.314696e-01    + i -5.555702e-01
		8'd25 : twiddle = { 16'd26790   , -16'd18868   }; //i=25 n=256 twiddle= 8.175848e-01    + i -5.758082e-01
		8'd26 : twiddle = { 16'd26319   , -16'd19519   }; //i=26 n=256 twiddle= 8.032075e-01    + i -5.956993e-01
		8'd27 : twiddle = { 16'd25832   , -16'd20159   }; //i=27 n=256 twiddle= 7.883464e-01    + i -6.152316e-01
		8'd28 : twiddle = { 16'd25329   , -16'd20787   }; //i=28 n=256 twiddle= 7.730105e-01    + i -6.343933e-01
		8'd29 : twiddle = { 16'd24811   , -16'd21403   }; //i=29 n=256 twiddle= 7.572088e-01    + i -6.531728e-01
		8'd30 : twiddle = { 16'd24279   , -16'd22005   }; //i=30 n=256 twiddle= 7.409511e-01    + i -6.715590e-01
		8'd31 : twiddle = { 16'd23731   , -16'd22594   }; //i=31 n=256 twiddle= 7.242471e-01    + i -6.895405e-01
		8'd32 : twiddle = { 16'd23170   , -16'd23170   }; //i=32 n=256 twiddle= 7.071068e-01    + i -7.071068e-01
		8'd33 : twiddle = { 16'd22594   , -16'd23731   }; //i=33 n=256 twiddle= 6.895405e-01    + i -7.242471e-01
		8'd34 : twiddle = { 16'd22005   , -16'd24279   }; //i=34 n=256 twiddle= 6.715590e-01    + i -7.409511e-01
		8'd35 : twiddle = { 16'd21403   , -16'd24811   }; //i=35 n=256 twiddle= 6.531728e-01    + i -7.572088e-01
		8'd36 : twiddle = { 16'd20787   , -16'd25329   }; //i=36 n=256 twiddle= 6.343933e-01    + i -7.730105e-01
		8'd37 : twiddle = { 16'd20159   , -16'd25832   }; //i=37 n=256 twiddle= 6.152316e-01    + i -7.883464e-01
		8'd38 : twiddle = { 16'd19519   , -16'd26319   }; //i=38 n=256 twiddle= 5.956993e-01    + i -8.032075e-01
		8'd39 : twiddle = { 16'd18868   , -16'd26790   }; //i=39 n=256 twiddle= 5.758082e-01    + i -8.175848e-01
		8'd40 : twiddle = { 16'd18204   , -16'd27245   }; //i=40 n=256 twiddle= 5.555702e-01    + i -8.314696e-01
		8'd41 : twiddle = { 16'd17530   , -16'd27683   }; //i=41 n=256 twiddle= 5.349976e-01    + i -8.448536e-01
		8'd42 : twiddle = { 16'd16846   , -16'd28105   }; //i=42 n=256 twiddle= 5.141027e-01    + i -8.577286e-01
		8'd43 : twiddle = { 16'd16151   , -16'd28510   }; //i=43 n=256 twiddle= 4.928982e-01    + i -8.700870e-01
		8'd44 : twiddle = { 16'd15446   , -16'd28898   }; //i=44 n=256 twiddle= 4.713967e-01    + i -8.819213e-01
		8'd45 : twiddle = { 16'd14732   , -16'd29268   }; //i=45 n=256 twiddle= 4.496113e-01    + i -8.932243e-01
		8'd46 : twiddle = { 16'd14010   , -16'd29621   }; //i=46 n=256 twiddle= 4.275551e-01    + i -9.039893e-01
		8'd47 : twiddle = { 16'd13279   , -16'd29956   }; //i=47 n=256 twiddle= 4.052413e-01    + i -9.142098e-01
		8'd48 : twiddle = { 16'd12539   , -16'd30273   }; //i=48 n=256 twiddle= 3.826834e-01    + i -9.238795e-01
		8'd49 : twiddle = { 16'd11793   , -16'd30571   }; //i=49 n=256 twiddle= 3.598950e-01    + i -9.329928e-01
		8'd50 : twiddle = { 16'd11039   , -16'd30852   }; //i=50 n=256 twiddle= 3.368899e-01    + i -9.415441e-01
		8'd51 : twiddle = { 16'd10278   , -16'd31113   }; //i=51 n=256 twiddle= 3.136817e-01    + i -9.495282e-01
		8'd52 : twiddle = { 16'd9512    , -16'd31356   }; //i=52 n=256 twiddle= 2.902847e-01    + i -9.569403e-01
		8'd53 : twiddle = { 16'd8739    , -16'd31580   }; //i=53 n=256 twiddle= 2.667128e-01    + i -9.637761e-01
		8'd54 : twiddle = { 16'd7962    , -16'd31785   }; //i=54 n=256 twiddle= 2.429802e-01    + i -9.700313e-01
		8'd55 : twiddle = { 16'd7179    , -16'd31971   }; //i=55 n=256 twiddle= 2.191012e-01    + i -9.757021e-01
		8'd56 : twiddle = { 16'd6393    , -16'd32137   }; //i=56 n=256 twiddle= 1.950903e-01    + i -9.807853e-01
		8'd57 : twiddle = { 16'd5602    , -16'd32285   }; //i=57 n=256 twiddle= 1.709619e-01    + i -9.852776e-01
		8'd58 : twiddle = { 16'd4808    , -16'd32412   }; //i=58 n=256 twiddle= 1.467305e-01    + i -9.891765e-01
		8'd59 : twiddle = { 16'd4011    , -16'd32521   }; //i=59 n=256 twiddle= 1.224107e-01    + i -9.924795e-01
		8'd60 : twiddle = { 16'd3212    , -16'd32609   }; //i=60 n=256 twiddle= 9.801714e-02    + i -9.951847e-01
		8'd61 : twiddle = { 16'd2410    , -16'd32678   }; //i=61 n=256 twiddle= 7.356456e-02    + i -9.972905e-01
		8'd62 : twiddle = { 16'd1608    , -16'd32728   }; //i=62 n=256 twiddle= 4.906767e-02    + i -9.987955e-01
		8'd63 : twiddle = { 16'd804     , -16'd32757   }; //i=63 n=256 twiddle= 2.454123e-02    + i -9.996988e-01
		8'd64 : twiddle = { 16'd0       , -16'd32767   }; //i=64 n=256 twiddle= 6.123234e-17    + i -1
		8'd65 : twiddle = {-16'd804     , -16'd32757   }; //i=65 n=256 twiddle= -2.454123e-02   + i -9.996988e-01
		8'd66 : twiddle = {-16'd1608    , -16'd32728   }; //i=66 n=256 twiddle= -4.906767e-02   + i -9.987955e-01
		8'd67 : twiddle = {-16'd2410    , -16'd32678   }; //i=67 n=256 twiddle= -7.356456e-02   + i -9.972905e-01
		8'd68 : twiddle = {-16'd3212    , -16'd32609   }; //i=68 n=256 twiddle= -9.801714e-02   + i -9.951847e-01
		8'd69 : twiddle = {-16'd4011    , -16'd32521   }; //i=69 n=256 twiddle= -1.224107e-01   + i -9.924795e-01
		8'd70 : twiddle = {-16'd4808    , -16'd32412   }; //i=70 n=256 twiddle= -1.467305e-01   + i -9.891765e-01
		8'd71 : twiddle = {-16'd5602    , -16'd32285   }; //i=71 n=256 twiddle= -1.709619e-01   + i -9.852776e-01
		8'd72 : twiddle = {-16'd6393    , -16'd32137   }; //i=72 n=256 twiddle= -1.950903e-01   + i -9.807853e-01
		8'd73 : twiddle = {-16'd7179    , -16'd31971   }; //i=73 n=256 twiddle= -2.191012e-01   + i -9.757021e-01
		8'd74 : twiddle = {-16'd7962    , -16'd31785   }; //i=74 n=256 twiddle= -2.429802e-01   + i -9.700313e-01
		8'd75 : twiddle = {-16'd8739    , -16'd31580   }; //i=75 n=256 twiddle= -2.667128e-01   + i -9.637761e-01
		8'd76 : twiddle = {-16'd9512    , -16'd31356   }; //i=76 n=256 twiddle= -2.902847e-01   + i -9.569403e-01
		8'd77 : twiddle = {-16'd10278   , -16'd31113   }; //i=77 n=256 twiddle= -3.136817e-01   + i -9.495282e-01
		8'd78 : twiddle = {-16'd11039   , -16'd30852   }; //i=78 n=256 twiddle= -3.368899e-01   + i -9.415441e-01
		8'd79 : twiddle = {-16'd11793   , -16'd30571   }; //i=79 n=256 twiddle= -3.598950e-01   + i -9.329928e-01
		8'd80 : twiddle = {-16'd12539   , -16'd30273   }; //i=80 n=256 twiddle= -3.826834e-01   + i -9.238795e-01
		8'd81 : twiddle = {-16'd13279   , -16'd29956   }; //i=81 n=256 twiddle= -4.052413e-01   + i -9.142098e-01
		8'd82 : twiddle = {-16'd14010   , -16'd29621   }; //i=82 n=256 twiddle= -4.275551e-01   + i -9.039893e-01
		8'd83 : twiddle = {-16'd14732   , -16'd29268   }; //i=83 n=256 twiddle= -4.496113e-01   + i -8.932243e-01
		8'd84 : twiddle = {-16'd15446   , -16'd28898   }; //i=84 n=256 twiddle= -4.713967e-01   + i -8.819213e-01
		8'd85 : twiddle = {-16'd16151   , -16'd28510   }; //i=85 n=256 twiddle= -4.928982e-01   + i -8.700870e-01
		8'd86 : twiddle = {-16'd16846   , -16'd28105   }; //i=86 n=256 twiddle= -5.141027e-01   + i -8.577286e-01
		8'd87 : twiddle = {-16'd17530   , -16'd27683   }; //i=87 n=256 twiddle= -5.349976e-01   + i -8.448536e-01
		8'd88 : twiddle = {-16'd18204   , -16'd27245   }; //i=88 n=256 twiddle= -5.555702e-01   + i -8.314696e-01
		8'd89 : twiddle = {-16'd18868   , -16'd26790   }; //i=89 n=256 twiddle= -5.758082e-01   + i -8.175848e-01
		8'd90 : twiddle = {-16'd19519   , -16'd26319   }; //i=90 n=256 twiddle= -5.956993e-01   + i -8.032075e-01
		8'd91 : twiddle = {-16'd20159   , -16'd25832   }; //i=91 n=256 twiddle= -6.152316e-01   + i -7.883464e-01
		8'd92 : twiddle = {-16'd20787   , -16'd25329   }; //i=92 n=256 twiddle= -6.343933e-01   + i -7.730105e-01
		8'd93 : twiddle = {-16'd21403   , -16'd24811   }; //i=93 n=256 twiddle= -6.531728e-01   + i -7.572088e-01
		8'd94 : twiddle = {-16'd22005   , -16'd24279   }; //i=94 n=256 twiddle= -6.715590e-01   + i -7.409511e-01
		8'd95 : twiddle = {-16'd22594   , -16'd23731   }; //i=95 n=256 twiddle= -6.895405e-01   + i -7.242471e-01
		8'd96 : twiddle = {-16'd23170   , -16'd23170   }; //i=96 n=256 twiddle= -7.071068e-01   + i -7.071068e-01
		8'd97 : twiddle = {-16'd23731   , -16'd22594   }; //i=97 n=256 twiddle= -7.242471e-01   + i -6.895405e-01
		8'd98 : twiddle = {-16'd24279   , -16'd22005   }; //i=98 n=256 twiddle= -7.409511e-01   + i -6.715590e-01
		8'd99 : twiddle = {-16'd24811   , -16'd21403   }; //i=99 n=256 twiddle= -7.572088e-01   + i -6.531728e-01
		8'd100: twiddle = {-16'd25329   , -16'd20787   }; //i=100 n=256 twiddle= -7.730105e-01   + i -6.343933e-01
		8'd101: twiddle = {-16'd25832   , -16'd20159   }; //i=101 n=256 twiddle= -7.883464e-01   + i -6.152316e-01
		8'd102: twiddle = {-16'd26319   , -16'd19519   }; //i=102 n=256 twiddle= -8.032075e-01   + i -5.956993e-01
		8'd103: twiddle = {-16'd26790   , -16'd18868   }; //i=103 n=256 twiddle= -8.175848e-01   + i -5.758082e-01
		8'd104: twiddle = {-16'd27245   , -16'd18204   }; //i=104 n=256 twiddle= -8.314696e-01   + i -5.555702e-01
		8'd105: twiddle = {-16'd27683   , -16'd17530   }; //i=105 n=256 twiddle= -8.448536e-01   + i -5.349976e-01
		8'd106: twiddle = {-16'd28105   , -16'd16846   }; //i=106 n=256 twiddle= -8.577286e-01   + i -5.141027e-01
		8'd107: twiddle = {-16'd28510   , -16'd16151   }; //i=107 n=256 twiddle= -8.700870e-01   + i -4.928982e-01
		8'd108: twiddle = {-16'd28898   , -16'd15446   }; //i=108 n=256 twiddle= -8.819213e-01   + i -4.713967e-01
		8'd109: twiddle = {-16'd29268   , -16'd14732   }; //i=109 n=256 twiddle= -8.932243e-01   + i -4.496113e-01
		8'd110: twiddle = {-16'd29621   , -16'd14010   }; //i=110 n=256 twiddle= -9.039893e-01   + i -4.275551e-01
		8'd111: twiddle = {-16'd29956   , -16'd13279   }; //i=111 n=256 twiddle= -9.142098e-01   + i -4.052413e-01
		8'd112: twiddle = {-16'd30273   , -16'd12539   }; //i=112 n=256 twiddle= -9.238795e-01   + i -3.826834e-01
		8'd113: twiddle = {-16'd30571   , -16'd11793   }; //i=113 n=256 twiddle= -9.329928e-01   + i -3.598950e-01
		8'd114: twiddle = {-16'd30852   , -16'd11039   }; //i=114 n=256 twiddle= -9.415441e-01   + i -3.368899e-01
		8'd115: twiddle = {-16'd31113   , -16'd10278   }; //i=115 n=256 twiddle= -9.495282e-01   + i -3.136817e-01
		8'd116: twiddle = {-16'd31356   , -16'd9512    }; //i=116 n=256 twiddle= -9.569403e-01   + i -2.902847e-01
		8'd117: twiddle = {-16'd31580   , -16'd8739    }; //i=117 n=256 twiddle= -9.637761e-01   + i -2.667128e-01
		8'd118: twiddle = {-16'd31785   , -16'd7962    }; //i=118 n=256 twiddle= -9.700313e-01   + i -2.429802e-01
		8'd119: twiddle = {-16'd31971   , -16'd7179    }; //i=119 n=256 twiddle= -9.757021e-01   + i -2.191012e-01
		8'd120: twiddle = {-16'd32137   , -16'd6393    }; //i=120 n=256 twiddle= -9.807853e-01   + i -1.950903e-01
		8'd121: twiddle = {-16'd32285   , -16'd5602    }; //i=121 n=256 twiddle= -9.852776e-01   + i -1.709619e-01
		8'd122: twiddle = {-16'd32412   , -16'd4808    }; //i=122 n=256 twiddle= -9.891765e-01   + i -1.467305e-01
		8'd123: twiddle = {-16'd32521   , -16'd4011    }; //i=123 n=256 twiddle= -9.924795e-01   + i -1.224107e-01
		8'd124: twiddle = {-16'd32609   , -16'd3212    }; //i=124 n=256 twiddle= -9.951847e-01   + i -9.801714e-02
		8'd125: twiddle = {-16'd32678   , -16'd2410    }; //i=125 n=256 twiddle= -9.972905e-01   + i -7.356456e-02
		8'd126: twiddle = {-16'd32728   , -16'd1608    }; //i=126 n=256 twiddle= -9.987955e-01   + i -4.906767e-02
		8'd127: twiddle = {-16'd32757   , -16'd804     }; //i=127 n=256 twiddle= -9.996988e-01   + i -2.454123e-02
		default: twiddle = 'bX;
		endcase
	end

endmodule