module HANN_LUT(n, hann);
	input [9:0] n;
		
	output reg [15:0] hann;
	
	always @ (n)
	begin
		//$display("LUT address=%d", n);
		case(n)
			10'd0  : hann = {16'd0       }; //i=0  n=1024 hann=    2.298488e-01
			10'd1  : hann = {16'd0       }; //i=1  n=1024 hann=    2.272723e-01
			10'd2  : hann = {16'd1       }; //i=2  n=1024 hann=    2.247061e-01
			10'd3  : hann = {16'd3       }; //i=3  n=1024 hann=    2.221503e-01
			10'd4  : hann = {16'd5       }; //i=4  n=1024 hann=    2.196048e-01
			10'd5  : hann = {16'd8       }; //i=5  n=1024 hann=    2.170700e-01
			10'd6  : hann = {16'd11      }; //i=6  n=1024 hann=    2.145458e-01
			10'd7  : hann = {16'd15      }; //i=7  n=1024 hann=    2.120324e-01
			10'd8  : hann = {16'd20      }; //i=8  n=1024 hann=    2.095297e-01
			10'd9  : hann = {16'd25      }; //i=9  n=1024 hann=    2.070381e-01
			10'd10 : hann = {16'd31      }; //i=10 n=1024 hann=    2.045574e-01
			10'd11 : hann = {16'd37      }; //i=11 n=1024 hann=    2.020879e-01
			10'd12 : hann = {16'd44      }; //i=12 n=1024 hann=    1.996296e-01
			10'd13 : hann = {16'd52      }; //i=13 n=1024 hann=    1.971826e-01
			10'd14 : hann = {16'd61      }; //i=14 n=1024 hann=    1.947470e-01
			10'd15 : hann = {16'd69      }; //i=15 n=1024 hann=    1.923229e-01
			10'd16 : hann = {16'd79      }; //i=16 n=1024 hann=    1.899104e-01
			10'd17 : hann = {16'd89      }; //i=17 n=1024 hann=    1.875096e-01
			10'd18 : hann = {16'd100     }; //i=18 n=1024 hann=    1.851205e-01
			10'd19 : hann = {16'd111     }; //i=19 n=1024 hann=    1.827433e-01
			10'd20 : hann = {16'd123     }; //i=20 n=1024 hann=    1.803780e-01
			10'd21 : hann = {16'd136     }; //i=21 n=1024 hann=    1.780248e-01
			10'd22 : hann = {16'd149     }; //i=22 n=1024 hann=    1.756836e-01
			10'd23 : hann = {16'd163     }; //i=23 n=1024 hann=    1.733547e-01
			10'd24 : hann = {16'd178     }; //i=24 n=1024 hann=    1.710381e-01
			10'd25 : hann = {16'd193     }; //i=25 n=1024 hann=    1.687339e-01
			10'd26 : hann = {16'd208     }; //i=26 n=1024 hann=    1.664421e-01
			10'd27 : hann = {16'd225     }; //i=27 n=1024 hann=    1.641629e-01
			10'd28 : hann = {16'd242     }; //i=28 n=1024 hann=    1.618964e-01
			10'd29 : hann = {16'd259     }; //i=29 n=1024 hann=    1.596426e-01
			10'd30 : hann = {16'd277     }; //i=30 n=1024 hann=    1.574015e-01
			10'd31 : hann = {16'd296     }; //i=31 n=1024 hann=    1.551734e-01
			10'd32 : hann = {16'd315     }; //i=32 n=1024 hann=    1.529583e-01
			10'd33 : hann = {16'd335     }; //i=33 n=1024 hann=    1.507562e-01
			10'd34 : hann = {16'd356     }; //i=34 n=1024 hann=    1.485673e-01
			10'd35 : hann = {16'd377     }; //i=35 n=1024 hann=    1.463916e-01
			10'd36 : hann = {16'd399     }; //i=36 n=1024 hann=    1.442293e-01
			10'd37 : hann = {16'd421     }; //i=37 n=1024 hann=    1.420803e-01
			10'd38 : hann = {16'd444     }; //i=38 n=1024 hann=    1.399448e-01
			10'd39 : hann = {16'd468     }; //i=39 n=1024 hann=    1.378229e-01
			10'd40 : hann = {16'd492     }; //i=40 n=1024 hann=    1.357146e-01
			10'd41 : hann = {16'd517     }; //i=41 n=1024 hann=    1.336200e-01
			10'd42 : hann = {16'd542     }; //i=42 n=1024 hann=    1.315392e-01
			10'd43 : hann = {16'd568     }; //i=43 n=1024 hann=    1.294722e-01
			10'd44 : hann = {16'd595     }; //i=44 n=1024 hann=    1.274193e-01
			10'd45 : hann = {16'd622     }; //i=45 n=1024 hann=    1.253803e-01
			10'd46 : hann = {16'd650     }; //i=46 n=1024 hann=    1.233555e-01
			10'd47 : hann = {16'd678     }; //i=47 n=1024 hann=    1.213448e-01
			10'd48 : hann = {16'd707     }; //i=48 n=1024 hann=    1.193484e-01
			10'd49 : hann = {16'd736     }; //i=49 n=1024 hann=    1.173663e-01
			10'd50 : hann = {16'd766     }; //i=50 n=1024 hann=    1.153987e-01
			10'd51 : hann = {16'd797     }; //i=51 n=1024 hann=    1.134455e-01
			10'd52 : hann = {16'd829     }; //i=52 n=1024 hann=    1.115068e-01
			10'd53 : hann = {16'd860     }; //i=53 n=1024 hann=    1.095828e-01
			10'd54 : hann = {16'd893     }; //i=54 n=1024 hann=    1.076735e-01
			10'd55 : hann = {16'd926     }; //i=55 n=1024 hann=    1.057790e-01
			10'd56 : hann = {16'd960     }; //i=56 n=1024 hann=    1.038993e-01
			10'd57 : hann = {16'd994     }; //i=57 n=1024 hann=    1.020345e-01
			10'd58 : hann = {16'd1029    }; //i=58 n=1024 hann=    1.001847e-01
			10'd59 : hann = {16'd1064    }; //i=59 n=1024 hann=    9.834993e-02
			10'd60 : hann = {16'd1100    }; //i=60 n=1024 hann=    9.653030e-02
			10'd61 : hann = {16'd1136    }; //i=61 n=1024 hann=    9.472587e-02
			10'd62 : hann = {16'd1174    }; //i=62 n=1024 hann=    9.293669e-02
			10'd63 : hann = {16'd1211    }; //i=63 n=1024 hann=    9.116284e-02
			10'd64 : hann = {16'd1250    }; //i=64 n=1024 hann=    8.940438e-02
			10'd65 : hann = {16'd1288    }; //i=65 n=1024 hann=    8.766138e-02
			10'd66 : hann = {16'd1328    }; //i=66 n=1024 hann=    8.593390e-02
			10'd67 : hann = {16'd1368    }; //i=67 n=1024 hann=    8.422201e-02
			10'd68 : hann = {16'd1408    }; //i=68 n=1024 hann=    8.252578e-02
			10'd69 : hann = {16'd1449    }; //i=69 n=1024 hann=    8.084526e-02
			10'd70 : hann = {16'd1491    }; //i=70 n=1024 hann=    7.918053e-02
			10'd71 : hann = {16'd1533    }; //i=71 n=1024 hann=    7.753163e-02
			10'd72 : hann = {16'd1576    }; //i=72 n=1024 hann=    7.589865e-02
			10'd73 : hann = {16'd1619    }; //i=73 n=1024 hann=    7.428163e-02
			10'd74 : hann = {16'd1663    }; //i=74 n=1024 hann=    7.268064e-02
			10'd75 : hann = {16'd1708    }; //i=75 n=1024 hann=    7.109574e-02
			10'd76 : hann = {16'd1753    }; //i=76 n=1024 hann=    6.952698e-02
			10'd77 : hann = {16'd1798    }; //i=77 n=1024 hann=    6.797443e-02
			10'd78 : hann = {16'd1844    }; //i=78 n=1024 hann=    6.643815e-02
			10'd79 : hann = {16'd1891    }; //i=79 n=1024 hann=    6.491819e-02
			10'd80 : hann = {16'd1938    }; //i=80 n=1024 hann=    6.341462e-02
			10'd81 : hann = {16'd1986    }; //i=81 n=1024 hann=    6.192747e-02
			10'd82 : hann = {16'd2034    }; //i=82 n=1024 hann=    6.045683e-02
			10'd83 : hann = {16'd2083    }; //i=83 n=1024 hann=    5.900273e-02
			10'd84 : hann = {16'd2133    }; //i=84 n=1024 hann=    5.756523e-02
			10'd85 : hann = {16'd2182    }; //i=85 n=1024 hann=    5.614439e-02
			10'd86 : hann = {16'd2233    }; //i=86 n=1024 hann=    5.474027e-02
			10'd87 : hann = {16'd2284    }; //i=87 n=1024 hann=    5.335290e-02
			10'd88 : hann = {16'd2335    }; //i=88 n=1024 hann=    5.198236e-02
			10'd89 : hann = {16'd2387    }; //i=89 n=1024 hann=    5.062868e-02
			10'd90 : hann = {16'd2440    }; //i=90 n=1024 hann=    4.929191e-02
			10'd91 : hann = {16'd2493    }; //i=91 n=1024 hann=    4.797212e-02
			10'd92 : hann = {16'd2547    }; //i=92 n=1024 hann=    4.666935e-02
			10'd93 : hann = {16'd2601    }; //i=93 n=1024 hann=    4.538364e-02
			10'd94 : hann = {16'd2655    }; //i=94 n=1024 hann=    4.411505e-02
			10'd95 : hann = {16'd2711    }; //i=95 n=1024 hann=    4.286363e-02
			10'd96 : hann = {16'd2766    }; //i=96 n=1024 hann=    4.162941e-02
			10'd97 : hann = {16'd2823    }; //i=97 n=1024 hann=    4.041245e-02
			10'd98 : hann = {16'd2879    }; //i=98 n=1024 hann=    3.921280e-02
			10'd99 : hann = {16'd2937    }; //i=99 n=1024 hann=    3.803049e-02
			10'd100: hann = {16'd2994    }; //i=100 n=1024 hann=    3.686558e-02
			10'd101: hann = {16'd3053    }; //i=101 n=1024 hann=    3.571810e-02
			10'd102: hann = {16'd3111    }; //i=102 n=1024 hann=    3.458810e-02
			10'd103: hann = {16'd3170    }; //i=103 n=1024 hann=    3.347563e-02
			10'd104: hann = {16'd3230    }; //i=104 n=1024 hann=    3.238072e-02
			10'd105: hann = {16'd3290    }; //i=105 n=1024 hann=    3.130341e-02
			10'd106: hann = {16'd3351    }; //i=106 n=1024 hann=    3.024376e-02
			10'd107: hann = {16'd3412    }; //i=107 n=1024 hann=    2.920178e-02
			10'd108: hann = {16'd3474    }; //i=108 n=1024 hann=    2.817754e-02
			10'd109: hann = {16'd3536    }; //i=109 n=1024 hann=    2.717105e-02
			10'd110: hann = {16'd3599    }; //i=110 n=1024 hann=    2.618237e-02
			10'd111: hann = {16'd3662    }; //i=111 n=1024 hann=    2.521153e-02
			10'd112: hann = {16'd3726    }; //i=112 n=1024 hann=    2.425856e-02
			10'd113: hann = {16'd3790    }; //i=113 n=1024 hann=    2.332351e-02
			10'd114: hann = {16'd3855    }; //i=114 n=1024 hann=    2.240640e-02
			10'd115: hann = {16'd3920    }; //i=115 n=1024 hann=    2.150727e-02
			10'd116: hann = {16'd3985    }; //i=116 n=1024 hann=    2.062616e-02
			10'd117: hann = {16'd4051    }; //i=117 n=1024 hann=    1.976309e-02
			10'd118: hann = {16'd4118    }; //i=118 n=1024 hann=    1.891811e-02
			10'd119: hann = {16'd4185    }; //i=119 n=1024 hann=    1.809124e-02
			10'd120: hann = {16'd4252    }; //i=120 n=1024 hann=    1.728251e-02
			10'd121: hann = {16'd4320    }; //i=121 n=1024 hann=    1.649196e-02
			10'd122: hann = {16'd4388    }; //i=122 n=1024 hann=    1.571961e-02
			10'd123: hann = {16'd4457    }; //i=123 n=1024 hann=    1.496549e-02
			10'd124: hann = {16'd4526    }; //i=124 n=1024 hann=    1.422963e-02
			10'd125: hann = {16'd4596    }; //i=125 n=1024 hann=    1.351207e-02
			10'd126: hann = {16'd4666    }; //i=126 n=1024 hann=    1.281282e-02
			10'd127: hann = {16'd4737    }; //i=127 n=1024 hann=    1.213191e-02
			10'd128: hann = {16'd4808    }; //i=128 n=1024 hann=    1.146937e-02
			10'd129: hann = {16'd4879    }; //i=129 n=1024 hann=    1.082522e-02
			10'd130: hann = {16'd4951    }; //i=130 n=1024 hann=    1.019949e-02
			10'd131: hann = {16'd5023    }; //i=131 n=1024 hann=    9.592200e-03
			10'd132: hann = {16'd5096    }; //i=132 n=1024 hann=    9.003374e-03
			10'd133: hann = {16'd5169    }; //i=133 n=1024 hann=    8.433033e-03
			10'd134: hann = {16'd5243    }; //i=134 n=1024 hann=    7.881200e-03
			10'd135: hann = {16'd5317    }; //i=135 n=1024 hann=    7.347895e-03
			10'd136: hann = {16'd5391    }; //i=136 n=1024 hann=    6.833138e-03
			10'd137: hann = {16'd5466    }; //i=137 n=1024 hann=    6.336948e-03
			10'd138: hann = {16'd5541    }; //i=138 n=1024 hann=    5.859344e-03
			10'd139: hann = {16'd5617    }; //i=139 n=1024 hann=    5.400345e-03
			10'd140: hann = {16'd5693    }; //i=140 n=1024 hann=    4.959967e-03
			10'd141: hann = {16'd5769    }; //i=141 n=1024 hann=    4.538226e-03
			10'd142: hann = {16'd5846    }; //i=142 n=1024 hann=    4.135140e-03
			10'd143: hann = {16'd5923    }; //i=143 n=1024 hann=    3.750723e-03
			10'd144: hann = {16'd6001    }; //i=144 n=1024 hann=    3.384989e-03
			10'd145: hann = {16'd6079    }; //i=145 n=1024 hann=    3.037953e-03
			10'd146: hann = {16'd6157    }; //i=146 n=1024 hann=    2.709627e-03
			10'd147: hann = {16'd6236    }; //i=147 n=1024 hann=    2.400023e-03
			10'd148: hann = {16'd6315    }; //i=148 n=1024 hann=    2.109154e-03
			10'd149: hann = {16'd6395    }; //i=149 n=1024 hann=    1.837030e-03
			10'd150: hann = {16'd6475    }; //i=150 n=1024 hann=    1.583662e-03
			10'd151: hann = {16'd6555    }; //i=151 n=1024 hann=    1.349059e-03
			10'd152: hann = {16'd6636    }; //i=152 n=1024 hann=    1.133230e-03
			10'd153: hann = {16'd6717    }; //i=153 n=1024 hann=    9.361827e-04
			10'd154: hann = {16'd6798    }; //i=154 n=1024 hann=    7.579250e-04
			10'd155: hann = {16'd6880    }; //i=155 n=1024 hann=    5.984636e-04
			10'd156: hann = {16'd6962    }; //i=156 n=1024 hann=    4.578043e-04
			10'd157: hann = {16'd7045    }; //i=157 n=1024 hann=    3.359525e-04
			10'd158: hann = {16'd7128    }; //i=158 n=1024 hann=    2.329127e-04
			10'd159: hann = {16'd7211    }; //i=159 n=1024 hann=    1.486889e-04
			10'd160: hann = {16'd7294    }; //i=160 n=1024 hann=    8.328426e-05
			10'd161: hann = {16'd7378    }; //i=161 n=1024 hann=    3.670117e-05
			10'd162: hann = {16'd7463    }; //i=162 n=1024 hann=    8.941417e-06
			10'd163: hann = {16'd7547    }; //i=163 n=1024 hann=    6.043018e-09
			10'd164: hann = {16'd7632    }; //i=164 n=1024 hann=    9.895386e-06
			10'd165: hann = {16'd7717    }; //i=165 n=1024 hann=    3.860907e-05
			10'd166: hann = {16'd7803    }; //i=166 n=1024 hann=    8.614603e-05
			10'd167: hann = {16'd7889    }; //i=167 n=1024 hann=    1.525045e-04
			10'd168: hann = {16'd7975    }; //i=168 n=1024 hann=    2.376819e-04
			10'd169: hann = {16'd8061    }; //i=169 n=1024 hann=    3.416750e-04
			10'd170: hann = {16'd8148    }; //i=170 n=1024 hann=    4.644800e-04
			10'd171: hann = {16'd8235    }; //i=171 n=1024 hann=    6.060923e-04
			10'd172: hann = {16'd8323    }; //i=172 n=1024 hann=    7.665065e-04
			10'd173: hann = {16'd8411    }; //i=173 n=1024 hann=    9.457165e-04
			10'd174: hann = {16'd8499    }; //i=174 n=1024 hann=    1.143716e-03
			10'd175: hann = {16'd8587    }; //i=175 n=1024 hann=    1.360496e-03
			10'd176: hann = {16'd8676    }; //i=176 n=1024 hann=    1.596051e-03
			10'd177: hann = {16'd8765    }; //i=177 n=1024 hann=    1.850370e-03
			10'd178: hann = {16'd8854    }; //i=178 n=1024 hann=    2.123443e-03
			10'd179: hann = {16'd8943    }; //i=179 n=1024 hann=    2.415262e-03
			10'd180: hann = {16'd9033    }; //i=180 n=1024 hann=    2.725815e-03
			10'd181: hann = {16'd9123    }; //i=181 n=1024 hann=    3.055089e-03
			10'd182: hann = {16'd9214    }; //i=182 n=1024 hann=    3.403074e-03
			10'd183: hann = {16'd9304    }; //i=183 n=1024 hann=    3.769755e-03
			10'd184: hann = {16'd9395    }; //i=184 n=1024 hann=    4.155118e-03
			10'd185: hann = {16'd9486    }; //i=185 n=1024 hann=    4.559150e-03
			10'd186: hann = {16'd9578    }; //i=186 n=1024 hann=    4.981835e-03
			10'd187: hann = {16'd9669    }; //i=187 n=1024 hann=    5.423157e-03
			10'd188: hann = {16'd9761    }; //i=188 n=1024 hann=    5.883100e-03
			10'd189: hann = {16'd9853    }; //i=189 n=1024 hann=    6.361646e-03
			10'd190: hann = {16'd9946    }; //i=190 n=1024 hann=    6.858777e-03
			10'd191: hann = {16'd10038   }; //i=191 n=1024 hann=    7.374475e-03
			10'd192: hann = {16'd10131   }; //i=192 n=1024 hann=    7.908720e-03
			10'd193: hann = {16'd10224   }; //i=193 n=1024 hann=    8.461491e-03
			10'd194: hann = {16'd10318   }; //i=194 n=1024 hann=    9.032769e-03
			10'd195: hann = {16'd10411   }; //i=195 n=1024 hann=    9.622531e-03
			10'd196: hann = {16'd10505   }; //i=196 n=1024 hann=    1.023076e-02
			10'd197: hann = {16'd10599   }; //i=197 n=1024 hann=    1.085742e-02
			10'd198: hann = {16'd10693   }; //i=198 n=1024 hann=    1.150250e-02
			10'd199: hann = {16'd10788   }; //i=199 n=1024 hann=    1.216597e-02
			10'd200: hann = {16'd10883   }; //i=200 n=1024 hann=    1.284781e-02
			10'd201: hann = {16'd10977   }; //i=201 n=1024 hann=    1.354799e-02
			10'd202: hann = {16'd11073   }; //i=202 n=1024 hann=    1.426649e-02
			10'd203: hann = {16'd11168   }; //i=203 n=1024 hann=    1.500327e-02
			10'd204: hann = {16'd11263   }; //i=204 n=1024 hann=    1.575831e-02
			10'd205: hann = {16'd11359   }; //i=205 n=1024 hann=    1.653158e-02
			10'd206: hann = {16'd11455   }; //i=206 n=1024 hann=    1.732306e-02
			10'd207: hann = {16'd11551   }; //i=207 n=1024 hann=    1.813271e-02
			10'd208: hann = {16'd11647   }; //i=208 n=1024 hann=    1.896050e-02
			10'd209: hann = {16'd11744   }; //i=209 n=1024 hann=    1.980640e-02
			10'd210: hann = {16'd11840   }; //i=210 n=1024 hann=    2.067038e-02
			10'd211: hann = {16'd11937   }; //i=211 n=1024 hann=    2.155240e-02
			10'd212: hann = {16'd12034   }; //i=212 n=1024 hann=    2.245244e-02
			10'd213: hann = {16'd12131   }; //i=213 n=1024 hann=    2.337046e-02
			10'd214: hann = {16'd12228   }; //i=214 n=1024 hann=    2.430643e-02
			10'd215: hann = {16'd12326   }; //i=215 n=1024 hann=    2.526030e-02
			10'd216: hann = {16'd12423   }; //i=216 n=1024 hann=    2.623205e-02
			10'd217: hann = {16'd12521   }; //i=217 n=1024 hann=    2.722163e-02
			10'd218: hann = {16'd12619   }; //i=218 n=1024 hann=    2.822902e-02
			10'd219: hann = {16'd12717   }; //i=219 n=1024 hann=    2.925416e-02
			10'd220: hann = {16'd12815   }; //i=220 n=1024 hann=    3.029703e-02
			10'd221: hann = {16'd12913   }; //i=221 n=1024 hann=    3.135758e-02
			10'd222: hann = {16'd13012   }; //i=222 n=1024 hann=    3.243578e-02
			10'd223: hann = {16'd13110   }; //i=223 n=1024 hann=    3.353158e-02
			10'd224: hann = {16'd13209   }; //i=224 n=1024 hann=    3.464495e-02
			10'd225: hann = {16'd13308   }; //i=225 n=1024 hann=    3.577583e-02
			10'd226: hann = {16'd13407   }; //i=226 n=1024 hann=    3.692419e-02
			10'd227: hann = {16'd13506   }; //i=227 n=1024 hann=    3.808999e-02
			10'd228: hann = {16'd13605   }; //i=228 n=1024 hann=    3.927317e-02
			10'd229: hann = {16'd13704   }; //i=229 n=1024 hann=    4.047371e-02
			10'd230: hann = {16'd13803   }; //i=230 n=1024 hann=    4.169154e-02
			10'd231: hann = {16'd13903   }; //i=231 n=1024 hann=    4.292663e-02
			10'd232: hann = {16'd14002   }; //i=232 n=1024 hann=    4.417893e-02
			10'd233: hann = {16'd14102   }; //i=233 n=1024 hann=    4.544839e-02
			10'd234: hann = {16'd14201   }; //i=234 n=1024 hann=    4.673496e-02
			10'd235: hann = {16'd14301   }; //i=235 n=1024 hann=    4.803860e-02
			10'd236: hann = {16'd14401   }; //i=236 n=1024 hann=    4.935925e-02
			10'd237: hann = {16'd14501   }; //i=237 n=1024 hann=    5.069687e-02
			10'd238: hann = {16'd14601   }; //i=238 n=1024 hann=    5.205141e-02
			10'd239: hann = {16'd14701   }; //i=239 n=1024 hann=    5.342281e-02
			10'd240: hann = {16'd14801   }; //i=240 n=1024 hann=    5.481102e-02
			10'd241: hann = {16'd14901   }; //i=241 n=1024 hann=    5.621600e-02
			10'd242: hann = {16'd15002   }; //i=242 n=1024 hann=    5.763768e-02
			10'd243: hann = {16'd15102   }; //i=243 n=1024 hann=    5.907602e-02
			10'd244: hann = {16'd15202   }; //i=244 n=1024 hann=    6.053096e-02
			10'd245: hann = {16'd15303   }; //i=245 n=1024 hann=    6.200244e-02
			10'd246: hann = {16'd15403   }; //i=246 n=1024 hann=    6.349042e-02
			10'd247: hann = {16'd15503   }; //i=247 n=1024 hann=    6.499483e-02
			10'd248: hann = {16'd15604   }; //i=248 n=1024 hann=    6.651561e-02
			10'd249: hann = {16'd15704   }; //i=249 n=1024 hann=    6.805272e-02
			10'd250: hann = {16'd15805   }; //i=250 n=1024 hann=    6.960609e-02
			10'd251: hann = {16'd15906   }; //i=251 n=1024 hann=    7.117566e-02
			10'd252: hann = {16'd16006   }; //i=252 n=1024 hann=    7.276138e-02
			10'd253: hann = {16'd16107   }; //i=253 n=1024 hann=    7.436319e-02
			10'd254: hann = {16'd16207   }; //i=254 n=1024 hann=    7.598102e-02
			10'd255: hann = {16'd16308   }; //i=255 n=1024 hann=    7.761481e-02
			10'd256: hann = {16'd16409   }; //i=256 n=1024 hann=    7.926451e-02
			10'd257: hann = {16'd16509   }; //i=257 n=1024 hann=    8.093004e-02
			10'd258: hann = {16'd16610   }; //i=258 n=1024 hann=    8.261136e-02
			10'd259: hann = {16'd16711   }; //i=259 n=1024 hann=    8.430839e-02
			10'd260: hann = {16'd16811   }; //i=260 n=1024 hann=    8.602107e-02
			10'd261: hann = {16'd16912   }; //i=261 n=1024 hann=    8.774933e-02
			10'd262: hann = {16'd17012   }; //i=262 n=1024 hann=    8.949312e-02
			10'd263: hann = {16'd17113   }; //i=263 n=1024 hann=    9.125236e-02
			10'd264: hann = {16'd17213   }; //i=264 n=1024 hann=    9.302699e-02
			10'd265: hann = {16'd17314   }; //i=265 n=1024 hann=    9.481694e-02
			10'd266: hann = {16'd17414   }; //i=266 n=1024 hann=    9.662215e-02
			10'd267: hann = {16'd17515   }; //i=267 n=1024 hann=    9.844255e-02
			10'd268: hann = {16'd17615   }; //i=268 n=1024 hann=    1.002781e-01
			10'd269: hann = {16'd17715   }; //i=269 n=1024 hann=    1.021286e-01
			10'd270: hann = {16'd17816   }; //i=270 n=1024 hann=    1.039942e-01
			10'd271: hann = {16'd17916   }; //i=271 n=1024 hann=    1.058746e-01
			10'd272: hann = {16'd18016   }; //i=272 n=1024 hann=    1.077699e-01
			10'd273: hann = {16'd18116   }; //i=273 n=1024 hann=    1.096800e-01
			10'd274: hann = {16'd18216   }; //i=274 n=1024 hann=    1.116047e-01
			10'd275: hann = {16'd18316   }; //i=275 n=1024 hann=    1.135441e-01
			10'd276: hann = {16'd18416   }; //i=276 n=1024 hann=    1.154980e-01
			10'd277: hann = {16'd18516   }; //i=277 n=1024 hann=    1.174664e-01
			10'd278: hann = {16'd18615   }; //i=278 n=1024 hann=    1.194492e-01
			10'd279: hann = {16'd18715   }; //i=279 n=1024 hann=    1.214464e-01
			10'd280: hann = {16'd18815   }; //i=280 n=1024 hann=    1.234577e-01
			10'd281: hann = {16'd18914   }; //i=281 n=1024 hann=    1.254833e-01
			10'd282: hann = {16'd19014   }; //i=282 n=1024 hann=    1.275230e-01
			10'd283: hann = {16'd19113   }; //i=283 n=1024 hann=    1.295766e-01
			10'd284: hann = {16'd19212   }; //i=284 n=1024 hann=    1.316443e-01
			10'd285: hann = {16'd19311   }; //i=285 n=1024 hann=    1.337258e-01
			10'd286: hann = {16'd19410   }; //i=286 n=1024 hann=    1.358211e-01
			10'd287: hann = {16'd19509   }; //i=287 n=1024 hann=    1.379301e-01
			10'd288: hann = {16'd19608   }; //i=288 n=1024 hann=    1.400527e-01
			10'd289: hann = {16'd19706   }; //i=289 n=1024 hann=    1.421889e-01
			10'd290: hann = {16'd19805   }; //i=290 n=1024 hann=    1.443385e-01
			10'd291: hann = {16'd19903   }; //i=291 n=1024 hann=    1.465016e-01
			10'd292: hann = {16'd20001   }; //i=292 n=1024 hann=    1.486779e-01
			10'd293: hann = {16'd20099   }; //i=293 n=1024 hann=    1.508675e-01
			10'd294: hann = {16'd20197   }; //i=294 n=1024 hann=    1.530702e-01
			10'd295: hann = {16'd20295   }; //i=295 n=1024 hann=    1.552860e-01
			10'd296: hann = {16'd20393   }; //i=296 n=1024 hann=    1.575148e-01
			10'd297: hann = {16'd20490   }; //i=297 n=1024 hann=    1.597565e-01
			10'd298: hann = {16'd20587   }; //i=298 n=1024 hann=    1.620109e-01
			10'd299: hann = {16'd20685   }; //i=299 n=1024 hann=    1.642781e-01
			10'd300: hann = {16'd20782   }; //i=300 n=1024 hann=    1.665580e-01
			10'd301: hann = {16'd20878   }; //i=301 n=1024 hann=    1.688504e-01
			10'd302: hann = {16'd20975   }; //i=302 n=1024 hann=    1.711552e-01
			10'd303: hann = {16'd21072   }; //i=303 n=1024 hann=    1.734724e-01
			10'd304: hann = {16'd21168   }; //i=304 n=1024 hann=    1.758020e-01
			10'd305: hann = {16'd21264   }; //i=305 n=1024 hann=    1.781437e-01
			10'd306: hann = {16'd21360   }; //i=306 n=1024 hann=    1.804976e-01
			10'd307: hann = {16'd21456   }; //i=307 n=1024 hann=    1.828635e-01
			10'd308: hann = {16'd21551   }; //i=308 n=1024 hann=    1.852413e-01
			10'd309: hann = {16'd21647   }; //i=309 n=1024 hann=    1.876310e-01
			10'd310: hann = {16'd21742   }; //i=310 n=1024 hann=    1.900324e-01
			10'd311: hann = {16'd21837   }; //i=311 n=1024 hann=    1.924455e-01
			10'd312: hann = {16'd21932   }; //i=312 n=1024 hann=    1.948702e-01
			10'd313: hann = {16'd22026   }; //i=313 n=1024 hann=    1.973063e-01
			10'd314: hann = {16'd22121   }; //i=314 n=1024 hann=    1.997539e-01
			10'd315: hann = {16'd22215   }; //i=315 n=1024 hann=    2.022128e-01
			10'd316: hann = {16'd22309   }; //i=316 n=1024 hann=    2.046829e-01
			10'd317: hann = {16'd22403   }; //i=317 n=1024 hann=    2.071641e-01
			10'd318: hann = {16'd22496   }; //i=318 n=1024 hann=    2.096563e-01
			10'd319: hann = {16'd22589   }; //i=319 n=1024 hann=    2.121595e-01
			10'd320: hann = {16'd22682   }; //i=320 n=1024 hann=    2.146735e-01
			10'd321: hann = {16'd22775   }; //i=321 n=1024 hann=    2.171982e-01
			10'd322: hann = {16'd22868   }; //i=322 n=1024 hann=    2.197336e-01
			10'd323: hann = {16'd22960   }; //i=323 n=1024 hann=    2.222795e-01
			10'd324: hann = {16'd23052   }; //i=324 n=1024 hann=    2.248359e-01
			10'd325: hann = {16'd23144   }; //i=325 n=1024 hann=    2.274027e-01
			10'd326: hann = {16'd23235   }; //i=326 n=1024 hann=    2.299797e-01
			10'd327: hann = {16'd23326   }; //i=327 n=1024 hann=    2.325669e-01
			10'd328: hann = {16'd23417   }; //i=328 n=1024 hann=    2.351641e-01
			10'd329: hann = {16'd23508   }; //i=329 n=1024 hann=    2.377713e-01
			10'd330: hann = {16'd23599   }; //i=330 n=1024 hann=    2.403884e-01
			10'd331: hann = {16'd23689   }; //i=331 n=1024 hann=    2.430153e-01
			10'd332: hann = {16'd23779   }; //i=332 n=1024 hann=    2.456519e-01
			10'd333: hann = {16'd23868   }; //i=333 n=1024 hann=    2.482980e-01
			10'd334: hann = {16'd23958   }; //i=334 n=1024 hann=    2.509536e-01
			10'd335: hann = {16'd24047   }; //i=335 n=1024 hann=    2.536185e-01
			10'd336: hann = {16'd24136   }; //i=336 n=1024 hann=    2.562928e-01
			10'd337: hann = {16'd24224   }; //i=337 n=1024 hann=    2.589762e-01
			10'd338: hann = {16'd24312   }; //i=338 n=1024 hann=    2.616687e-01
			10'd339: hann = {16'd24400   }; //i=339 n=1024 hann=    2.643702e-01
			10'd340: hann = {16'd24488   }; //i=340 n=1024 hann=    2.670805e-01
			10'd341: hann = {16'd24575   }; //i=341 n=1024 hann=    2.697996e-01
			10'd342: hann = {16'd24662   }; //i=342 n=1024 hann=    2.725274e-01
			10'd343: hann = {16'd24749   }; //i=343 n=1024 hann=    2.752638e-01
			10'd344: hann = {16'd24835   }; //i=344 n=1024 hann=    2.780086e-01
			10'd345: hann = {16'd24921   }; //i=345 n=1024 hann=    2.807617e-01
			10'd346: hann = {16'd25007   }; //i=346 n=1024 hann=    2.835232e-01
			10'd347: hann = {16'd25092   }; //i=347 n=1024 hann=    2.862927e-01
			10'd348: hann = {16'd25178   }; //i=348 n=1024 hann=    2.890703e-01
			10'd349: hann = {16'd25262   }; //i=349 n=1024 hann=    2.918559e-01
			10'd350: hann = {16'd25347   }; //i=350 n=1024 hann=    2.946493e-01
			10'd351: hann = {16'd25431   }; //i=351 n=1024 hann=    2.974504e-01
			10'd352: hann = {16'd25514   }; //i=352 n=1024 hann=    3.002592e-01
			10'd353: hann = {16'd25598   }; //i=353 n=1024 hann=    3.030754e-01
			10'd354: hann = {16'd25681   }; //i=354 n=1024 hann=    3.058991e-01
			10'd355: hann = {16'd25764   }; //i=355 n=1024 hann=    3.087301e-01
			10'd356: hann = {16'd25846   }; //i=356 n=1024 hann=    3.115683e-01
			10'd357: hann = {16'd25928   }; //i=357 n=1024 hann=    3.144136e-01
			10'd358: hann = {16'd26009   }; //i=358 n=1024 hann=    3.172659e-01
			10'd359: hann = {16'd26091   }; //i=359 n=1024 hann=    3.201250e-01
			10'd360: hann = {16'd26172   }; //i=360 n=1024 hann=    3.229909e-01
			10'd361: hann = {16'd26252   }; //i=361 n=1024 hann=    3.258635e-01
			10'd362: hann = {16'd26332   }; //i=362 n=1024 hann=    3.287427e-01
			10'd363: hann = {16'd26412   }; //i=363 n=1024 hann=    3.316283e-01
			10'd364: hann = {16'd26491   }; //i=364 n=1024 hann=    3.345202e-01
			10'd365: hann = {16'd26570   }; //i=365 n=1024 hann=    3.374184e-01
			10'd366: hann = {16'd26649   }; //i=366 n=1024 hann=    3.403226e-01
			10'd367: hann = {16'd26727   }; //i=367 n=1024 hann=    3.432329e-01
			10'd368: hann = {16'd26805   }; //i=368 n=1024 hann=    3.461491e-01
			10'd369: hann = {16'd26882   }; //i=369 n=1024 hann=    3.490711e-01
			10'd370: hann = {16'd26960   }; //i=370 n=1024 hann=    3.519988e-01
			10'd371: hann = {16'd27036   }; //i=371 n=1024 hann=    3.549321e-01
			10'd372: hann = {16'd27112   }; //i=372 n=1024 hann=    3.578708e-01
			10'd373: hann = {16'd27188   }; //i=373 n=1024 hann=    3.608148e-01
			10'd374: hann = {16'd27264   }; //i=374 n=1024 hann=    3.637641e-01
			10'd375: hann = {16'd27339   }; //i=375 n=1024 hann=    3.667185e-01
			10'd376: hann = {16'd27413   }; //i=376 n=1024 hann=    3.696780e-01
			10'd377: hann = {16'd27488   }; //i=377 n=1024 hann=    3.726423e-01
			10'd378: hann = {16'd27561   }; //i=378 n=1024 hann=    3.756115e-01
			10'd379: hann = {16'd27635   }; //i=379 n=1024 hann=    3.785853e-01
			10'd380: hann = {16'd27708   }; //i=380 n=1024 hann=    3.815637e-01
			10'd381: hann = {16'd27780   }; //i=381 n=1024 hann=    3.845466e-01
			10'd382: hann = {16'd27852   }; //i=382 n=1024 hann=    3.875338e-01
			10'd383: hann = {16'd27924   }; //i=383 n=1024 hann=    3.905252e-01
			10'd384: hann = {16'd27995   }; //i=384 n=1024 hann=    3.935208e-01
			10'd385: hann = {16'd28066   }; //i=385 n=1024 hann=    3.965204e-01
			10'd386: hann = {16'd28136   }; //i=386 n=1024 hann=    3.995238e-01
			10'd387: hann = {16'd28206   }; //i=387 n=1024 hann=    4.025311e-01
			10'd388: hann = {16'd28275   }; //i=388 n=1024 hann=    4.055420e-01
			10'd389: hann = {16'd28344   }; //i=389 n=1024 hann=    4.085565e-01
			10'd390: hann = {16'd28413   }; //i=390 n=1024 hann=    4.115744e-01
			10'd391: hann = {16'd28481   }; //i=391 n=1024 hann=    4.145956e-01
			10'd392: hann = {16'd28549   }; //i=392 n=1024 hann=    4.176201e-01
			10'd393: hann = {16'd28616   }; //i=393 n=1024 hann=    4.206477e-01
			10'd394: hann = {16'd28683   }; //i=394 n=1024 hann=    4.236782e-01
			10'd395: hann = {16'd28749   }; //i=395 n=1024 hann=    4.267117e-01
			10'd396: hann = {16'd28815   }; //i=396 n=1024 hann=    4.297478e-01
			10'd397: hann = {16'd28880   }; //i=397 n=1024 hann=    4.327867e-01
			10'd398: hann = {16'd28945   }; //i=398 n=1024 hann=    4.358280e-01
			10'd399: hann = {16'd29009   }; //i=399 n=1024 hann=    4.388718e-01
			10'd400: hann = {16'd29073   }; //i=400 n=1024 hann=    4.419179e-01
			10'd401: hann = {16'd29136   }; //i=401 n=1024 hann=    4.449662e-01
			10'd402: hann = {16'd29199   }; //i=402 n=1024 hann=    4.480165e-01
			10'd403: hann = {16'd29262   }; //i=403 n=1024 hann=    4.510688e-01
			10'd404: hann = {16'd29324   }; //i=404 n=1024 hann=    4.541229e-01
			10'd405: hann = {16'd29385   }; //i=405 n=1024 hann=    4.571788e-01
			10'd406: hann = {16'd29446   }; //i=406 n=1024 hann=    4.602363e-01
			10'd407: hann = {16'd29507   }; //i=407 n=1024 hann=    4.632952e-01
			10'd408: hann = {16'd29567   }; //i=408 n=1024 hann=    4.663556e-01
			10'd409: hann = {16'd29626   }; //i=409 n=1024 hann=    4.694172e-01
			10'd410: hann = {16'd29685   }; //i=410 n=1024 hann=    4.724800e-01
			10'd411: hann = {16'd29744   }; //i=411 n=1024 hann=    4.755438e-01
			10'd412: hann = {16'd29802   }; //i=412 n=1024 hann=    4.786085e-01
			10'd413: hann = {16'd29859   }; //i=413 n=1024 hann=    4.816741e-01
			10'd414: hann = {16'd29916   }; //i=414 n=1024 hann=    4.847403e-01
			10'd415: hann = {16'd29973   }; //i=415 n=1024 hann=    4.878071e-01
			10'd416: hann = {16'd30029   }; //i=416 n=1024 hann=    4.908744e-01
			10'd417: hann = {16'd30084   }; //i=417 n=1024 hann=    4.939420e-01
			10'd418: hann = {16'd30139   }; //i=418 n=1024 hann=    4.970098e-01
			10'd419: hann = {16'd30193   }; //i=419 n=1024 hann=    5.000777e-01
			10'd420: hann = {16'd30247   }; //i=420 n=1024 hann=    5.031457e-01
			10'd421: hann = {16'd30301   }; //i=421 n=1024 hann=    5.062135e-01
			10'd422: hann = {16'd30353   }; //i=422 n=1024 hann=    5.092811e-01
			10'd423: hann = {16'd30406   }; //i=423 n=1024 hann=    5.123483e-01
			10'd424: hann = {16'd30457   }; //i=424 n=1024 hann=    5.154151e-01
			10'd425: hann = {16'd30509   }; //i=425 n=1024 hann=    5.184813e-01
			10'd426: hann = {16'd30559   }; //i=426 n=1024 hann=    5.215468e-01
			10'd427: hann = {16'd30610   }; //i=427 n=1024 hann=    5.246115e-01
			10'd428: hann = {16'd30659   }; //i=428 n=1024 hann=    5.276752e-01
			10'd429: hann = {16'd30708   }; //i=429 n=1024 hann=    5.307380e-01
			10'd430: hann = {16'd30757   }; //i=430 n=1024 hann=    5.337995e-01
			10'd431: hann = {16'd30805   }; //i=431 n=1024 hann=    5.368598e-01
			10'd432: hann = {16'd30852   }; //i=432 n=1024 hann=    5.399187e-01
			10'd433: hann = {16'd30899   }; //i=433 n=1024 hann=    5.429761e-01
			10'd434: hann = {16'd30946   }; //i=434 n=1024 hann=    5.460319e-01
			10'd435: hann = {16'd30992   }; //i=435 n=1024 hann=    5.490859e-01
			10'd436: hann = {16'd31037   }; //i=436 n=1024 hann=    5.521381e-01
			10'd437: hann = {16'd31082   }; //i=437 n=1024 hann=    5.551884e-01
			10'd438: hann = {16'd31126   }; //i=438 n=1024 hann=    5.582365e-01
			10'd439: hann = {16'd31169   }; //i=439 n=1024 hann=    5.612825e-01
			10'd440: hann = {16'd31212   }; //i=440 n=1024 hann=    5.643261e-01
			10'd441: hann = {16'd31255   }; //i=441 n=1024 hann=    5.673674e-01
			10'd442: hann = {16'd31297   }; //i=442 n=1024 hann=    5.704061e-01
			10'd443: hann = {16'd31338   }; //i=443 n=1024 hann=    5.734421e-01
			10'd444: hann = {16'd31379   }; //i=444 n=1024 hann=    5.764754e-01
			10'd445: hann = {16'd31419   }; //i=445 n=1024 hann=    5.795058e-01
			10'd446: hann = {16'd31459   }; //i=446 n=1024 hann=    5.825332e-01
			10'd447: hann = {16'd31498   }; //i=447 n=1024 hann=    5.855575e-01
			10'd448: hann = {16'd31537   }; //i=448 n=1024 hann=    5.885786e-01
			10'd449: hann = {16'd31575   }; //i=449 n=1024 hann=    5.915964e-01
			10'd450: hann = {16'd31612   }; //i=450 n=1024 hann=    5.946107e-01
			10'd451: hann = {16'd31649   }; //i=451 n=1024 hann=    5.976214e-01
			10'd452: hann = {16'd31685   }; //i=452 n=1024 hann=    6.006285e-01
			10'd453: hann = {16'd31721   }; //i=453 n=1024 hann=    6.036317e-01
			10'd454: hann = {16'd31756   }; //i=454 n=1024 hann=    6.066311e-01
			10'd455: hann = {16'd31790   }; //i=455 n=1024 hann=    6.096265e-01
			10'd456: hann = {16'd31824   }; //i=456 n=1024 hann=    6.126177e-01
			10'd457: hann = {16'd31858   }; //i=457 n=1024 hann=    6.156047e-01
			10'd458: hann = {16'd31890   }; //i=458 n=1024 hann=    6.185873e-01
			10'd459: hann = {16'd31923   }; //i=459 n=1024 hann=    6.215655e-01
			10'd460: hann = {16'd31954   }; //i=460 n=1024 hann=    6.245391e-01
			10'd461: hann = {16'd31985   }; //i=461 n=1024 hann=    6.275080e-01
			10'd462: hann = {16'd32016   }; //i=462 n=1024 hann=    6.304721e-01
			10'd463: hann = {16'd32045   }; //i=463 n=1024 hann=    6.334313e-01
			10'd464: hann = {16'd32075   }; //i=464 n=1024 hann=    6.363855e-01
			10'd465: hann = {16'd32103   }; //i=465 n=1024 hann=    6.393345e-01
			10'd466: hann = {16'd32131   }; //i=466 n=1024 hann=    6.422783e-01
			10'd467: hann = {16'd32159   }; //i=467 n=1024 hann=    6.452167e-01
			10'd468: hann = {16'd32186   }; //i=468 n=1024 hann=    6.481497e-01
			10'd469: hann = {16'd32212   }; //i=469 n=1024 hann=    6.510771e-01
			10'd470: hann = {16'd32238   }; //i=470 n=1024 hann=    6.539988e-01
			10'd471: hann = {16'd32263   }; //i=471 n=1024 hann=    6.569147e-01
			10'd472: hann = {16'd32287   }; //i=472 n=1024 hann=    6.598247e-01
			10'd473: hann = {16'd32311   }; //i=473 n=1024 hann=    6.627287e-01
			10'd474: hann = {16'd32334   }; //i=474 n=1024 hann=    6.656265e-01
			10'd475: hann = {16'd32357   }; //i=475 n=1024 hann=    6.685181e-01
			10'd476: hann = {16'd32379   }; //i=476 n=1024 hann=    6.714034e-01
			10'd477: hann = {16'd32401   }; //i=477 n=1024 hann=    6.742822e-01
			10'd478: hann = {16'd32421   }; //i=478 n=1024 hann=    6.771545e-01
			10'd479: hann = {16'd32442   }; //i=479 n=1024 hann=    6.800200e-01
			10'd480: hann = {16'd32461   }; //i=480 n=1024 hann=    6.828789e-01
			10'd481: hann = {16'd32480   }; //i=481 n=1024 hann=    6.857308e-01
			10'd482: hann = {16'd32499   }; //i=482 n=1024 hann=    6.885757e-01
			10'd483: hann = {16'd32517   }; //i=483 n=1024 hann=    6.914135e-01
			10'd484: hann = {16'd32534   }; //i=484 n=1024 hann=    6.942442e-01
			10'd485: hann = {16'd32550   }; //i=485 n=1024 hann=    6.970675e-01
			10'd486: hann = {16'd32566   }; //i=486 n=1024 hann=    6.998834e-01
			10'd487: hann = {16'd32582   }; //i=487 n=1024 hann=    7.026917e-01
			10'd488: hann = {16'd32597   }; //i=488 n=1024 hann=    7.054925e-01
			10'd489: hann = {16'd32611   }; //i=489 n=1024 hann=    7.082855e-01
			10'd490: hann = {16'd32624   }; //i=490 n=1024 hann=    7.110706e-01
			10'd491: hann = {16'd32637   }; //i=491 n=1024 hann=    7.138478e-01
			10'd492: hann = {16'd32650   }; //i=492 n=1024 hann=    7.166170e-01
			10'd493: hann = {16'd32661   }; //i=493 n=1024 hann=    7.193780e-01
			10'd494: hann = {16'd32672   }; //i=494 n=1024 hann=    7.221307e-01
			10'd495: hann = {16'd32683   }; //i=495 n=1024 hann=    7.248751e-01
			10'd496: hann = {16'd32693   }; //i=496 n=1024 hann=    7.276110e-01
			10'd497: hann = {16'd32702   }; //i=497 n=1024 hann=    7.303384e-01
			10'd498: hann = {16'd32711   }; //i=498 n=1024 hann=    7.330570e-01
			10'd499: hann = {16'd32719   }; //i=499 n=1024 hann=    7.357669e-01
			10'd500: hann = {16'd32726   }; //i=500 n=1024 hann=    7.384679e-01
			10'd501: hann = {16'd32733   }; //i=501 n=1024 hann=    7.411600e-01
			10'd502: hann = {16'd32739   }; //i=502 n=1024 hann=    7.438429e-01
			10'd503: hann = {16'd32745   }; //i=503 n=1024 hann=    7.465167e-01
			10'd504: hann = {16'd32750   }; //i=504 n=1024 hann=    7.491812e-01
			10'd505: hann = {16'd32754   }; //i=505 n=1024 hann=    7.518364e-01
			10'd506: hann = {16'd32758   }; //i=506 n=1024 hann=    7.544820e-01
			10'd507: hann = {16'd32761   }; //i=507 n=1024 hann=    7.571180e-01
			10'd508: hann = {16'd32763   }; //i=508 n=1024 hann=    7.597444e-01
			10'd509: hann = {16'd32765   }; //i=509 n=1024 hann=    7.623610e-01
			10'd510: hann = {16'd32766   }; //i=510 n=1024 hann=    7.649677e-01
			10'd511: hann = {16'd32767   }; //i=511 n=1024 hann=    7.675645e-01
			default: hann = 'bX;
		endcase
	end

endmodule