`timescale 1ns / 1ps

module FFT1024_tb_v;
	parameter PRE = 16;
		
	reg Clk;
	reg Reset, Start;
	reg signed [PRE-1:0] X_Re [1024:0];
	reg signed [PRE-1:0] X_Im [1024:0];
	
	// Outputs
	wire signed [2*PRE-1:0] X_Re_out [1024:0];
	wire signed [2*PRE-1:0] X_Im_out [1024:0];
	wire Done;
	
	// Instantiate the Unit Under Test (UUT)
	FFT1024 uut (
		.Clk(Clk),
		.Reset(Reset),
		.Start(Start),
		.x_re(X_Re[PRE-1:0]),
		.x_im(X_Im),
		.Done(Done)
	);
	
	
	initial
	begin
		Clk = 0; // Initialize clock
		Start = 0;
		Reset = 0;
	end
	
	// Keep clock running
	always
	begin
		#20; 
		Clk = ~ Clk; 
	end
	
	initial
	begin
		Start = 0;
		#200
		// FFT
		X_Re[0] = 15'd87845;
		X_Re[1] = 15'd3344;
		X_Re[2] = 15'd8055;
		X_Re[3] = -15'd3237;
		X_Re[4] = -15'd3178;
		X_Re[5] = -15'd8097;
		X_Re[6] = -15'd13493;
		X_Re[7] = -15'd45742;
		X_Re[8] = -15'd5662;
		X_Re[9] = -15'd166613;
		X_Re[10] = -15'd45666;
		X_Re[11] = 15'd71943;
		X_Re[12] = -15'd7187;
		X_Re[13] = -15'd40016;
		X_Re[14] = 15'd2080;
		X_Re[15] = 15'd16013;
		X_Re[16] = -15'd12426;
		X_Re[17] = 15'd41019;
		X_Re[18] = -15'd32079;
		X_Re[19] = -15'd54871;
		X_Re[20] = 15'd1037;
		X_Re[21] = -15'd19342;
		X_Re[22] = -15'd4748;
		X_Re[23] = 15'd13800;
		X_Re[24] = -15'd5577;
		X_Re[25] = 15'd2592;
		X_Re[26] = 15'd41646;
		X_Re[27] = -15'd73347;
		X_Re[28] = -15'd34797;
		X_Re[29] = -15'd23890;
		X_Re[30] = -15'd38433;
		X_Re[31] = -15'd23713;
		X_Re[32] = -15'd20014;
		X_Re[33] = -15'd10798;
		X_Re[34] = -15'd22086;
		X_Re[35] = 15'd31774;
		X_Re[36] = -15'd57943;
		X_Re[37] = -15'd33674;
		X_Re[38] = -15'd92155;
		X_Re[39] = -15'd219111;
		X_Re[40] = 15'd422815;
		X_Re[41] = 15'd77266;
		X_Re[42] = 15'd48085;
		X_Re[43] = 15'd19080;
		X_Re[44] = 15'd71278;
		X_Re[45] = 15'd32371;
		X_Re[46] = 15'd7926;
		X_Re[47] = 15'd35091;
		X_Re[48] = 15'd37484;
		X_Re[49] = 15'd19509;
		X_Re[50] = 15'd18707;
		X_Re[51] = 15'd44296;
		X_Re[52] = 15'd3041;
		X_Re[53] = 15'd200812;
		X_Re[54] = -15'd32042;
		X_Re[55] = -15'd2465;
		X_Re[56] = 15'd19028;
		X_Re[57] = 15'd16164;
		X_Re[58] = 15'd99801;
		X_Re[59] = 15'd172680;
		X_Re[60] = -15'd374488;
		X_Re[61] = -15'd76563;
		X_Re[62] = -15'd68355;
		X_Re[63] = -15'd73725;
		X_Re[64] = -15'd89550;
		X_Re[65] = -15'd84078;
		X_Re[66] = -15'd350559;
		X_Re[67] = -15'd220475;
		X_Re[68] = 15'd25897;
		X_Re[69] = 15'd98286;
		X_Re[70] = 15'd24689;
		X_Re[71] = 15'd86424;
		X_Re[72] = 15'd20529;
		X_Re[73] = 15'd27560;
		X_Re[74] = 15'd24094;
		X_Re[75] = 15'd20953;
		X_Re[76] = 15'd15514;
		X_Re[77] = 15'd18835;
		X_Re[78] = -15'd2159;
		X_Re[79] = -15'd322659;
		X_Re[80] = -15'd103143;
		X_Re[81] = 15'd21865;
		X_Re[82] = 15'd5014;
		X_Re[83] = 15'd10478;
		X_Re[84] = 15'd7487;
		X_Re[85] = 15'd1599;
		X_Re[86] = 15'd508;
		X_Re[87] = 15'd6553;
		X_Re[88] = 15'd12647;
		X_Re[89] = 15'd328;
		X_Re[90] = 15'd13322;
		X_Re[91] = 15'd19519;
		X_Re[92] = 15'd10361;
		X_Re[93] = 15'd11635;
		X_Re[94] = 15'd53368;
		X_Re[95] = -15'd32083;
		X_Re[96] = -15'd1423;
		X_Re[97] = -15'd15483;
		X_Re[98] = -15'd6194;
		X_Re[99] = 15'd3784;
		X_Re[100] = 15'd2743;
		X_Re[101] = 15'd2850;
		X_Re[102] = -15'd429;
		X_Re[103] = -15'd6999;
		X_Re[104] = -15'd8783;
		X_Re[105] = -15'd33732;
		X_Re[106] = 15'd36890;
		X_Re[107] = 15'd20766;
		X_Re[108] = 15'd2968;
		X_Re[109] = 15'd13462;
		X_Re[110] = -15'd870;
		X_Re[111] = 15'd7264;
		X_Re[112] = -15'd4449;
		X_Re[113] = 15'd4331;
		X_Re[114] = 15'd8206;
		X_Re[115] = 15'd3472;
		X_Re[116] = 15'd7848;
		X_Re[117] = 15'd24008;
		X_Re[118] = -15'd14034;
		X_Re[119] = -15'd93185;
		X_Re[120] = 15'd35868;
		X_Re[121] = -15'd8956;
		X_Re[122] = 15'd16199;
		X_Re[123] = 15'd4346;
		X_Re[124] = -15'd653;
		X_Re[125] = 15'd11710;
		X_Re[126] = 15'd242;
		X_Re[127] = -15'd2025;
		X_Re[128] = -15'd2026;
		X_Re[129] = -15'd5956;
		X_Re[130] = 15'd1626;
		X_Re[131] = -15'd5217;
		X_Re[132] = 15'd28921;
		X_Re[133] = 15'd348596;
		X_Re[134] = 15'd70108;
		X_Re[135] = -15'd59599;
		X_Re[136] = 15'd4423;
		X_Re[137] = -15'd10221;
		X_Re[138] = -15'd2938;
		X_Re[139] = -15'd7719;
		X_Re[140] = -15'd14770;
		X_Re[141] = 15'd24684;
		X_Re[142] = 15'd8862;
		X_Re[143] = -15'd7572;
		X_Re[144] = 15'd2346;
		X_Re[145] = 15'd1621;
		X_Re[146] = 15'd7001;
		X_Re[147] = 15'd5648;
		X_Re[148] = 15'd1191;
		X_Re[149] = 15'd3541;
		X_Re[150] = 15'd8099;
		X_Re[151] = 15'd9251;
		X_Re[152] = 15'd4481;
		X_Re[153] = 15'd5927;
		X_Re[154] = -15'd785;
		X_Re[155] = 15'd7908;
		X_Re[156] = -15'd9583;
		X_Re[157] = 15'd16551;
		X_Re[158] = 15'd43192;
		X_Re[159] = -15'd26098;
		X_Re[160] = 15'd44207;
		X_Re[161] = -15'd53731;
		X_Re[162] = -15'd13945;
		X_Re[163] = 15'd7595;
		X_Re[164] = -15'd18047;
		X_Re[165] = -15'd7142;
		X_Re[166] = 15'd2843;
		X_Re[167] = -15'd9092;
		X_Re[168] = -15'd5662;
		X_Re[169] = 15'd6326;
		X_Re[170] = -15'd4492;
		X_Re[171] = -15'd4310;
		X_Re[172] = -15'd6699;
		X_Re[173] = 15'd3645;
		X_Re[174] = -15'd5322;
		X_Re[175] = 15'd72;
		X_Re[176] = -15'd8022;
		X_Re[177] = -15'd10941;
		X_Re[178] = 15'd21188;
		X_Re[179] = -15'd36128;
		X_Re[180] = 15'd6839;
		X_Re[181] = 15'd7248;
		X_Re[182] = -15'd1081;
		X_Re[183] = -15'd10342;
		X_Re[184] = -15'd5390;
		X_Re[185] = -15'd1703;
		X_Re[186] = -15'd9567;
		X_Re[187] = -15'd2829;
		X_Re[188] = -15'd1650;
		X_Re[189] = 15'd33592;
		X_Re[190] = -15'd5174;
		X_Re[191] = -15'd4157;
		X_Re[192] = -15'd4998;
		X_Re[193] = -15'd13655;
		X_Re[194] = -15'd12119;
		X_Re[195] = -15'd25781;
		X_Re[196] = -15'd36556;
		X_Re[197] = -15'd22939;
		X_Re[198] = 15'd11030;
		X_Re[199] = 15'd73677;
		X_Re[200] = 15'd79471;
		X_Re[201] = -15'd12893;
		X_Re[202] = 15'd45500;
		X_Re[203] = 15'd22040;
		X_Re[204] = 15'd113;
		X_Re[205] = 15'd14818;
		X_Re[206] = 15'd13157;
		X_Re[207] = 15'd8849;
		X_Re[208] = 15'd7302;
		X_Re[209] = 15'd3742;
		X_Re[210] = 15'd1597;
		X_Re[211] = -15'd4435;
		X_Re[212] = 15'd12250;
		X_Re[213] = 15'd14568;
		X_Re[214] = 15'd5259;
		X_Re[215] = 15'd6701;
		X_Re[216] = 15'd1389;
		X_Re[217] = 15'd5842;
		X_Re[218] = 15'd4029;
		X_Re[219] = -15'd4858;
		X_Re[220] = -15'd3645;
		X_Re[221] = -15'd672;
		X_Re[222] = 15'd4974;
		X_Re[223] = 15'd18305;
		X_Re[224] = 15'd1586;
		X_Re[225] = 15'd3644;
		X_Re[226] = -15'd3440;
		X_Re[227] = -15'd1443;
		X_Re[228] = 15'd2725;
		X_Re[229] = -15'd1024;
		X_Re[230] = 15'd5750;
		X_Re[231] = 15'd2656;
		X_Re[232] = -15'd1000;
		X_Re[233] = -15'd3814;
		X_Re[234] = 15'd12974;
		X_Re[235] = 15'd444;
		X_Re[236] = -15'd135;
		X_Re[237] = -15'd17114;
		X_Re[238] = -15'd20408;
		X_Re[239] = 15'd15575;
		X_Re[240] = 15'd23887;
		X_Re[241] = -15'd5678;
		X_Re[242] = 15'd2716;
		X_Re[243] = 15'd7430;
		X_Re[244] = 15'd5149;
		X_Re[245] = 15'd1347;
		X_Re[246] = 15'd198;
		X_Re[247] = 15'd4325;
		X_Re[248] = 15'd1647;
		X_Re[249] = 15'd2362;
		X_Re[250] = -15'd4211;
		X_Re[251] = -15'd4557;
		X_Re[252] = 15'd247;
		X_Re[253] = 15'd561;
		X_Re[254] = -15'd2300;
		X_Re[255] = -15'd2812;
		X_Re[256] = 15'd4199;
		X_Re[257] = 15'd6102;
		X_Re[258] = 15'd2286;
		X_Re[259] = -15'd1321;
		X_Re[260] = 15'd3711;
		X_Re[261] = -15'd4232;
		X_Re[262] = -15'd1814;
		X_Re[263] = -15'd1966;
		X_Re[264] = -15'd20260;
		X_Re[265] = -15'd12043;
		X_Re[266] = -15'd27418;
		X_Re[267] = 15'd74501;
		X_Re[268] = -15'd12580;
		X_Re[269] = 15'd51561;
		X_Re[270] = 15'd38212;
		X_Re[271] = 15'd5018;
		X_Re[272] = 15'd10433;
		X_Re[273] = 15'd1041;
		X_Re[274] = 15'd4839;
		X_Re[275] = -15'd2275;
		X_Re[276] = 15'd1240;
		X_Re[277] = -15'd9718;
		X_Re[278] = 15'd19251;
		X_Re[279] = 15'd15875;
		X_Re[280] = 15'd24907;
		X_Re[281] = -15'd17830;
		X_Re[282] = 15'd22972;
		X_Re[283] = -15'd15060;
		X_Re[284] = -15'd17454;
		X_Re[285] = 15'd14979;
		X_Re[286] = 15'd5478;
		X_Re[287] = 15'd8163;
		X_Re[288] = 15'd9653;
		X_Re[289] = 15'd7815;
		X_Re[290] = -15'd4390;
		X_Re[291] = -15'd1107;
		X_Re[292] = 15'd4921;
		X_Re[293] = 15'd5641;
		X_Re[294] = 15'd8048;
		X_Re[295] = 15'd20142;
		X_Re[296] = 15'd304;
		X_Re[297] = -15'd21717;
		X_Re[298] = -15'd15387;
		X_Re[299] = 15'd910;
		X_Re[300] = -15'd5584;
		X_Re[301] = -15'd2360;
		X_Re[302] = -15'd4573;
		X_Re[303] = 15'd4507;
		X_Re[304] = -15'd468;
		X_Re[305] = -15'd2353;
		X_Re[306] = -15'd4686;
		X_Re[307] = -15'd997;
		X_Re[308] = 15'd3014;
		X_Re[309] = -15'd3343;
		X_Re[310] = -15'd10076;
		X_Re[311] = -15'd4711;
		X_Re[312] = -15'd119;
		X_Re[313] = -15'd8284;
		X_Re[314] = -15'd6385;
		X_Re[315] = 15'd1001;
		X_Re[316] = -15'd20754;
		X_Re[317] = 15'd6510;
		X_Re[318] = 15'd9622;
		X_Re[319] = -15'd12026;
		X_Re[320] = 15'd2135;
		X_Re[321] = 15'd4892;
		X_Re[322] = 15'd14113;
		X_Re[323] = 15'd12783;
		X_Re[324] = 15'd9026;
		X_Re[325] = -15'd3351;
		X_Re[326] = -15'd3522;
		X_Re[327] = -15'd1883;
		X_Re[328] = -15'd2104;
		X_Re[329] = 15'd2955;
		X_Re[330] = 15'd1624;
		X_Re[331] = 15'd9906;
		X_Re[332] = -15'd31088;
		X_Re[333] = -15'd69284;
		X_Re[334] = -15'd21741;
		X_Re[335] = 15'd26174;
		X_Re[336] = 15'd21107;
		X_Re[337] = 15'd27095;
		X_Re[338] = 15'd17744;
		X_Re[339] = 15'd7843;
		X_Re[340] = 15'd3575;
		X_Re[341] = 15'd5268;
		X_Re[342] = 15'd2275;
		X_Re[343] = 15'd5093;
		X_Re[344] = 15'd4152;
		X_Re[345] = 15'd6587;
		X_Re[346] = 15'd5706;
		X_Re[347] = 15'd9694;
		X_Re[348] = -15'd219;
		X_Re[349] = -15'd6394;
		X_Re[350] = 15'd9541;
		X_Re[351] = 15'd419;
		X_Re[352] = -15'd6571;
		X_Re[353] = -15'd12040;
		X_Re[354] = 15'd12326;
		X_Re[355] = 15'd13884;
		X_Re[356] = -15'd2894;
		X_Re[357] = 15'd10079;
		X_Re[358] = 15'd498;
		X_Re[359] = -15'd3106;
		X_Re[360] = 15'd11603;
		X_Re[361] = -15'd2867;
		X_Re[362] = 15'd3477;
		X_Re[363] = -15'd5876;
		X_Re[364] = -15'd3806;
		X_Re[365] = -15'd14665;
		X_Re[366] = 15'd4292;
		X_Re[367] = 15'd2298;
		X_Re[368] = 15'd1134;
		X_Re[369] = 15'd4562;
		X_Re[370] = -15'd4028;
		X_Re[371] = 15'd1076;
		X_Re[372] = 15'd1307;
		X_Re[373] = 15'd1266;
		X_Re[374] = 15'd5262;
		X_Re[375] = -15'd3120;
		X_Re[376] = 15'd2932;
		X_Re[377] = 15'd1223;
		X_Re[378] = 15'd4195;
		X_Re[379] = 15'd8723;
		X_Re[380] = 15'd2828;
		X_Re[381] = -15'd2569;
		X_Re[382] = 15'd185;
		X_Re[383] = 15'd791;
		X_Re[384] = 15'd3287;
		X_Re[385] = 15'd2779;
		X_Re[386] = 15'd1264;
		X_Re[387] = 15'd1993;
		X_Re[388] = -15'd2303;
		X_Re[389] = -15'd5224;
		X_Re[390] = 15'd4668;
		X_Re[391] = -15'd484;
		X_Re[392] = -15'd1336;
		X_Re[393] = 15'd3668;
		X_Re[394] = 15'd7126;
		X_Re[395] = -15'd696;
		X_Re[396] = 15'd5664;
		X_Re[397] = 15'd6114;
		X_Re[398] = 15'd5014;
		X_Re[399] = -15'd6974;
		X_Re[400] = 15'd6777;
		X_Re[401] = -15'd5889;
		X_Re[402] = 15'd8449;
		X_Re[403] = -15'd10760;
		X_Re[404] = -15'd14396;
		X_Re[405] = 15'd3588;
		X_Re[406] = -15'd2938;
		X_Re[407] = 15'd1930;
		X_Re[408] = 15'd524;
		X_Re[409] = -15'd10544;
		X_Re[410] = -15'd1736;
		X_Re[411] = -15'd11328;
		X_Re[412] = 15'd1017;
		X_Re[413] = -15'd2833;
		X_Re[414] = -15'd6321;
		X_Re[415] = -15'd7040;
		X_Re[416] = -15'd1046;
		X_Re[417] = -15'd4148;
		X_Re[418] = 15'd8989;
		X_Re[419] = 15'd14251;
		X_Re[420] = 15'd1665;
		X_Re[421] = 15'd9134;
		X_Re[422] = -15'd3527;
		X_Re[423] = 15'd487;
		X_Re[424] = -15'd8390;
		X_Re[425] = -15'd7080;
		X_Re[426] = -15'd1364;
		X_Re[427] = -15'd5337;
		X_Re[428] = -15'd3161;
		X_Re[429] = 15'd4474;
		X_Re[430] = 15'd771;
		X_Re[431] = 15'd11294;
		X_Re[432] = 15'd710;
		X_Re[433] = 15'd4136;
		X_Re[434] = -15'd1406;
		X_Re[435] = 15'd1701;
		X_Re[436] = 15'd3648;
		X_Re[437] = -15'd2515;
		X_Re[438] = 15'd5600;
		X_Re[439] = -15'd1077;
		X_Re[440] = -15'd5290;
		X_Re[441] = -15'd1696;
		X_Re[442] = 15'd253;
		X_Re[443] = -15'd3289;
		X_Re[444] = -15'd3339;
		X_Re[445] = 15'd2039;
		X_Re[446] = -15'd239;
		X_Re[447] = -15'd744;
		X_Re[448] = -15'd438;
		X_Re[449] = -15'd648;
		X_Re[450] = 15'd4640;
		X_Re[451] = -15'd785;
		X_Re[452] = 15'd3136;
		X_Re[453] = -15'd1347;
		X_Re[454] = -15'd2142;
		X_Re[455] = 15'd81;
		X_Re[456] = -15'd610;
		X_Re[457] = 15'd3765;
		X_Re[458] = 15'd4386;
		X_Re[459] = 15'd5782;
		X_Re[460] = -15'd4289;
		X_Re[461] = -15'd2578;
		X_Re[462] = -15'd7178;
		X_Re[463] = 15'd2181;
		X_Re[464] = -15'd983;
		X_Re[465] = 15'd478;
		X_Re[466] = -15'd12519;
		X_Re[467] = -15'd5800;
		X_Re[468] = -15'd11525;
		X_Re[469] = -15'd3360;
		X_Re[470] = -15'd9081;
		X_Re[471] = -15'd5005;
		X_Re[472] = 15'd12347;
		X_Re[473] = 15'd6589;
		X_Re[474] = -15'd4590;
		X_Re[475] = -15'd7421;
		X_Re[476] = -15'd7911;
		X_Re[477] = -15'd3481;
		X_Re[478] = 15'd503;
		X_Re[479] = -15'd4816;
		X_Re[480] = -15'd66;
		X_Re[481] = -15'd3201;
		X_Re[482] = -15'd4789;
		X_Re[483] = 15'd468;
		X_Re[484] = 15'd259;
		X_Re[485] = 15'd2268;
		X_Re[486] = 15'd14370;
		X_Re[487] = 15'd7708;
		X_Re[488] = 15'd12342;
		X_Re[489] = -15'd582;
		X_Re[490] = 15'd3663;
		X_Re[491] = -15'd3903;
		X_Re[492] = -15'd8920;
		X_Re[493] = -15'd857;
		X_Re[494] = -15'd4053;
		X_Re[495] = -15'd1268;
		X_Re[496] = 15'd5599;
		X_Re[497] = 15'd3546;
		X_Re[498] = -15'd1949;
		X_Re[499] = -15'd2754;
		X_Re[500] = 15'd5736;
		X_Re[501] = 15'd725;
		X_Re[502] = -15'd6801;
		X_Re[503] = 15'd4936;
		X_Re[504] = -15'd1656;
		X_Re[505] = -15'd1849;
		X_Re[506] = -15'd7295;
		X_Re[507] = 15'd7049;
		X_Re[508] = -15'd804;
		X_Re[509] = 15'd3487;
		X_Re[510] = -15'd2807;
		X_Re[511] = 15'd1575;
		X_Re[512] = -15'd1627;
		X_Re[513] = 15'd1575;
		X_Re[514] = -15'd2807;
		X_Re[515] = 15'd3487;
		X_Re[516] = -15'd804;
		X_Re[517] = 15'd7049;
		X_Re[518] = -15'd7295;
		X_Re[519] = -15'd1849;
		X_Re[520] = -15'd1656;
		X_Re[521] = 15'd4936;
		X_Re[522] = -15'd6801;
		X_Re[523] = 15'd725;
		X_Re[524] = 15'd5736;
		X_Re[525] = -15'd2754;
		X_Re[526] = -15'd1949;
		X_Re[527] = 15'd3546;
		X_Re[528] = 15'd5599;
		X_Re[529] = -15'd1268;
		X_Re[530] = -15'd4053;
		X_Re[531] = -15'd857;
		X_Re[532] = -15'd8920;
		X_Re[533] = -15'd3903;
		X_Re[534] = 15'd3663;
		X_Re[535] = -15'd582;
		X_Re[536] = 15'd12342;
		X_Re[537] = 15'd7708;
		X_Re[538] = 15'd14370;
		X_Re[539] = 15'd2268;
		X_Re[540] = 15'd259;
		X_Re[541] = 15'd468;
		X_Re[542] = -15'd4789;
		X_Re[543] = -15'd3201;
		X_Re[544] = -15'd66;
		X_Re[545] = -15'd4816;
		X_Re[546] = 15'd503;
		X_Re[547] = -15'd3481;
		X_Re[548] = -15'd7911;
		X_Re[549] = -15'd7421;
		X_Re[550] = -15'd4590;
		X_Re[551] = 15'd6589;
		X_Re[552] = 15'd12347;
		X_Re[553] = -15'd5005;
		X_Re[554] = -15'd9081;
		X_Re[555] = -15'd3360;
		X_Re[556] = -15'd11525;
		X_Re[557] = -15'd5800;
		X_Re[558] = -15'd12519;
		X_Re[559] = 15'd478;
		X_Re[560] = -15'd983;
		X_Re[561] = 15'd2181;
		X_Re[562] = -15'd7178;
		X_Re[563] = -15'd2578;
		X_Re[564] = -15'd4289;
		X_Re[565] = 15'd5782;
		X_Re[566] = 15'd4386;
		X_Re[567] = 15'd3765;
		X_Re[568] = -15'd610;
		X_Re[569] = 15'd81;
		X_Re[570] = -15'd2142;
		X_Re[571] = -15'd1347;
		X_Re[572] = 15'd3136;
		X_Re[573] = -15'd785;
		X_Re[574] = 15'd4640;
		X_Re[575] = -15'd648;
		X_Re[576] = -15'd438;
		X_Re[577] = -15'd744;
		X_Re[578] = -15'd239;
		X_Re[579] = 15'd2039;
		X_Re[580] = -15'd3339;
		X_Re[581] = -15'd3289;
		X_Re[582] = 15'd253;
		X_Re[583] = -15'd1696;
		X_Re[584] = -15'd5290;
		X_Re[585] = -15'd1077;
		X_Re[586] = 15'd5600;
		X_Re[587] = -15'd2515;
		X_Re[588] = 15'd3648;
		X_Re[589] = 15'd1701;
		X_Re[590] = -15'd1406;
		X_Re[591] = 15'd4136;
		X_Re[592] = 15'd710;
		X_Re[593] = 15'd11294;
		X_Re[594] = 15'd771;
		X_Re[595] = 15'd4474;
		X_Re[596] = -15'd3161;
		X_Re[597] = -15'd5337;
		X_Re[598] = -15'd1364;
		X_Re[599] = -15'd7080;
		X_Re[600] = -15'd8390;
		X_Re[601] = 15'd487;
		X_Re[602] = -15'd3527;
		X_Re[603] = 15'd9134;
		X_Re[604] = 15'd1665;
		X_Re[605] = 15'd14251;
		X_Re[606] = 15'd8989;
		X_Re[607] = -15'd4148;
		X_Re[608] = -15'd1046;
		X_Re[609] = -15'd7040;
		X_Re[610] = -15'd6321;
		X_Re[611] = -15'd2833;
		X_Re[612] = 15'd1017;
		X_Re[613] = -15'd11328;
		X_Re[614] = -15'd1736;
		X_Re[615] = -15'd10544;
		X_Re[616] = 15'd524;
		X_Re[617] = 15'd1930;
		X_Re[618] = -15'd2938;
		X_Re[619] = 15'd3588;
		X_Re[620] = -15'd14396;
		X_Re[621] = -15'd10760;
		X_Re[622] = 15'd8449;
		X_Re[623] = -15'd5889;
		X_Re[624] = 15'd6777;
		X_Re[625] = -15'd6974;
		X_Re[626] = 15'd5014;
		X_Re[627] = 15'd6114;
		X_Re[628] = 15'd5664;
		X_Re[629] = -15'd696;
		X_Re[630] = 15'd7126;
		X_Re[631] = 15'd3668;
		X_Re[632] = -15'd1336;
		X_Re[633] = -15'd484;
		X_Re[634] = 15'd4668;
		X_Re[635] = -15'd5224;
		X_Re[636] = -15'd2303;
		X_Re[637] = 15'd1993;
		X_Re[638] = 15'd1264;
		X_Re[639] = 15'd2779;
		X_Re[640] = 15'd3287;
		X_Re[641] = 15'd791;
		X_Re[642] = 15'd185;
		X_Re[643] = -15'd2569;
		X_Re[644] = 15'd2828;
		X_Re[645] = 15'd8723;
		X_Re[646] = 15'd4195;
		X_Re[647] = 15'd1223;
		X_Re[648] = 15'd2932;
		X_Re[649] = -15'd3120;
		X_Re[650] = 15'd5262;
		X_Re[651] = 15'd1266;
		X_Re[652] = 15'd1307;
		X_Re[653] = 15'd1076;
		X_Re[654] = -15'd4028;
		X_Re[655] = 15'd4562;
		X_Re[656] = 15'd1134;
		X_Re[657] = 15'd2298;
		X_Re[658] = 15'd4292;
		X_Re[659] = -15'd14665;
		X_Re[660] = -15'd3806;
		X_Re[661] = -15'd5876;
		X_Re[662] = 15'd3477;
		X_Re[663] = -15'd2867;
		X_Re[664] = 15'd11603;
		X_Re[665] = -15'd3106;
		X_Re[666] = 15'd498;
		X_Re[667] = 15'd10079;
		X_Re[668] = -15'd2894;
		X_Re[669] = 15'd13884;
		X_Re[670] = 15'd12326;
		X_Re[671] = -15'd12040;
		X_Re[672] = -15'd6571;
		X_Re[673] = 15'd419;
		X_Re[674] = 15'd9541;
		X_Re[675] = -15'd6394;
		X_Re[676] = -15'd219;
		X_Re[677] = 15'd9694;
		X_Re[678] = 15'd5706;
		X_Re[679] = 15'd6587;
		X_Re[680] = 15'd4152;
		X_Re[681] = 15'd5093;
		X_Re[682] = 15'd2275;
		X_Re[683] = 15'd5268;
		X_Re[684] = 15'd3575;
		X_Re[685] = 15'd7843;
		X_Re[686] = 15'd17744;
		X_Re[687] = 15'd27095;
		X_Re[688] = 15'd21107;
		X_Re[689] = 15'd26174;
		X_Re[690] = -15'd21741;
		X_Re[691] = -15'd69284;
		X_Re[692] = -15'd31088;
		X_Re[693] = 15'd9906;
		X_Re[694] = 15'd1624;
		X_Re[695] = 15'd2955;
		X_Re[696] = -15'd2104;
		X_Re[697] = -15'd1883;
		X_Re[698] = -15'd3522;
		X_Re[699] = -15'd3351;
		X_Re[700] = 15'd9026;
		X_Re[701] = 15'd12783;
		X_Re[702] = 15'd14113;
		X_Re[703] = 15'd4892;
		X_Re[704] = 15'd2135;
		X_Re[705] = -15'd12026;
		X_Re[706] = 15'd9622;
		X_Re[707] = 15'd6510;
		X_Re[708] = -15'd20754;
		X_Re[709] = 15'd1001;
		X_Re[710] = -15'd6385;
		X_Re[711] = -15'd8284;
		X_Re[712] = -15'd119;
		X_Re[713] = -15'd4711;
		X_Re[714] = -15'd10076;
		X_Re[715] = -15'd3343;
		X_Re[716] = 15'd3014;
		X_Re[717] = -15'd997;
		X_Re[718] = -15'd4686;
		X_Re[719] = -15'd2353;
		X_Re[720] = -15'd468;
		X_Re[721] = 15'd4507;
		X_Re[722] = -15'd4573;
		X_Re[723] = -15'd2360;
		X_Re[724] = -15'd5584;
		X_Re[725] = 15'd910;
		X_Re[726] = -15'd15387;
		X_Re[727] = -15'd21717;
		X_Re[728] = 15'd304;
		X_Re[729] = 15'd20142;
		X_Re[730] = 15'd8048;
		X_Re[731] = 15'd5641;
		X_Re[732] = 15'd4921;
		X_Re[733] = -15'd1107;
		X_Re[734] = -15'd4390;
		X_Re[735] = 15'd7815;
		X_Re[736] = 15'd9653;
		X_Re[737] = 15'd8163;
		X_Re[738] = 15'd5478;
		X_Re[739] = 15'd14979;
		X_Re[740] = -15'd17454;
		X_Re[741] = -15'd15060;
		X_Re[742] = 15'd22972;
		X_Re[743] = -15'd17830;
		X_Re[744] = 15'd24907;
		X_Re[745] = 15'd15875;
		X_Re[746] = 15'd19251;
		X_Re[747] = -15'd9718;
		X_Re[748] = 15'd1240;
		X_Re[749] = -15'd2275;
		X_Re[750] = 15'd4839;
		X_Re[751] = 15'd1041;
		X_Re[752] = 15'd10433;
		X_Re[753] = 15'd5018;
		X_Re[754] = 15'd38212;
		X_Re[755] = 15'd51561;
		X_Re[756] = -15'd12580;
		X_Re[757] = 15'd74501;
		X_Re[758] = -15'd27418;
		X_Re[759] = -15'd12043;
		X_Re[760] = -15'd20260;
		X_Re[761] = -15'd1966;
		X_Re[762] = -15'd1814;
		X_Re[763] = -15'd4232;
		X_Re[764] = 15'd3711;
		X_Re[765] = -15'd1321;
		X_Re[766] = 15'd2286;
		X_Re[767] = 15'd6102;
		X_Re[768] = 15'd4199;
		X_Re[769] = -15'd2812;
		X_Re[770] = -15'd2300;
		X_Re[771] = 15'd561;
		X_Re[772] = 15'd247;
		X_Re[773] = -15'd4557;
		X_Re[774] = -15'd4211;
		X_Re[775] = 15'd2362;
		X_Re[776] = 15'd1647;
		X_Re[777] = 15'd4325;
		X_Re[778] = 15'd198;
		X_Re[779] = 15'd1347;
		X_Re[780] = 15'd5149;
		X_Re[781] = 15'd7430;
		X_Re[782] = 15'd2716;
		X_Re[783] = -15'd5678;
		X_Re[784] = 15'd23887;
		X_Re[785] = 15'd15575;
		X_Re[786] = -15'd20408;
		X_Re[787] = -15'd17114;
		X_Re[788] = -15'd135;
		X_Re[789] = 15'd444;
		X_Re[790] = 15'd12974;
		X_Re[791] = -15'd3814;
		X_Re[792] = -15'd1000;
		X_Re[793] = 15'd2656;
		X_Re[794] = 15'd5750;
		X_Re[795] = -15'd1024;
		X_Re[796] = 15'd2725;
		X_Re[797] = -15'd1443;
		X_Re[798] = -15'd3440;
		X_Re[799] = 15'd3644;
		X_Re[800] = 15'd1586;
		X_Re[801] = 15'd18305;
		X_Re[802] = 15'd4974;
		X_Re[803] = -15'd672;
		X_Re[804] = -15'd3645;
		X_Re[805] = -15'd4858;
		X_Re[806] = 15'd4029;
		X_Re[807] = 15'd5842;
		X_Re[808] = 15'd1389;
		X_Re[809] = 15'd6701;
		X_Re[810] = 15'd5259;
		X_Re[811] = 15'd14568;
		X_Re[812] = 15'd12250;
		X_Re[813] = -15'd4435;
		X_Re[814] = 15'd1597;
		X_Re[815] = 15'd3742;
		X_Re[816] = 15'd7302;
		X_Re[817] = 15'd8849;
		X_Re[818] = 15'd13157;
		X_Re[819] = 15'd14818;
		X_Re[820] = 15'd113;
		X_Re[821] = 15'd22040;
		X_Re[822] = 15'd45500;
		X_Re[823] = -15'd12893;
		X_Re[824] = 15'd79471;
		X_Re[825] = 15'd73677;
		X_Re[826] = 15'd11030;
		X_Re[827] = -15'd22939;
		X_Re[828] = -15'd36556;
		X_Re[829] = -15'd25781;
		X_Re[830] = -15'd12119;
		X_Re[831] = -15'd13655;
		X_Re[832] = -15'd4998;
		X_Re[833] = -15'd4157;
		X_Re[834] = -15'd5174;
		X_Re[835] = 15'd33592;
		X_Re[836] = -15'd1650;
		X_Re[837] = -15'd2829;
		X_Re[838] = -15'd9567;
		X_Re[839] = -15'd1703;
		X_Re[840] = -15'd5390;
		X_Re[841] = -15'd10342;
		X_Re[842] = -15'd1081;
		X_Re[843] = 15'd7248;
		X_Re[844] = 15'd6839;
		X_Re[845] = -15'd36128;
		X_Re[846] = 15'd21188;
		X_Re[847] = -15'd10941;
		X_Re[848] = -15'd8022;
		X_Re[849] = 15'd72;
		X_Re[850] = -15'd5322;
		X_Re[851] = 15'd3645;
		X_Re[852] = -15'd6699;
		X_Re[853] = -15'd4310;
		X_Re[854] = -15'd4492;
		X_Re[855] = 15'd6326;
		X_Re[856] = -15'd5662;
		X_Re[857] = -15'd9092;
		X_Re[858] = 15'd2843;
		X_Re[859] = -15'd7142;
		X_Re[860] = -15'd18047;
		X_Re[861] = 15'd7595;
		X_Re[862] = -15'd13945;
		X_Re[863] = -15'd53731;
		X_Re[864] = 15'd44207;
		X_Re[865] = -15'd26098;
		X_Re[866] = 15'd43192;
		X_Re[867] = 15'd16551;
		X_Re[868] = -15'd9583;
		X_Re[869] = 15'd7908;
		X_Re[870] = -15'd785;
		X_Re[871] = 15'd5927;
		X_Re[872] = 15'd4481;
		X_Re[873] = 15'd9251;
		X_Re[874] = 15'd8099;
		X_Re[875] = 15'd3541;
		X_Re[876] = 15'd1191;
		X_Re[877] = 15'd5648;
		X_Re[878] = 15'd7001;
		X_Re[879] = 15'd1621;
		X_Re[880] = 15'd2346;
		X_Re[881] = -15'd7572;
		X_Re[882] = 15'd8862;
		X_Re[883] = 15'd24684;
		X_Re[884] = -15'd14770;
		X_Re[885] = -15'd7719;
		X_Re[886] = -15'd2938;
		X_Re[887] = -15'd10221;
		X_Re[888] = 15'd4423;
		X_Re[889] = -15'd59599;
		X_Re[890] = 15'd70108;
		X_Re[891] = 15'd348596;
		X_Re[892] = 15'd28921;
		X_Re[893] = -15'd5217;
		X_Re[894] = 15'd1626;
		X_Re[895] = -15'd5956;
		X_Re[896] = -15'd2026;
		X_Re[897] = -15'd2025;
		X_Re[898] = 15'd242;
		X_Re[899] = 15'd11710;
		X_Re[900] = -15'd653;
		X_Re[901] = 15'd4346;
		X_Re[902] = 15'd16199;
		X_Re[903] = -15'd8956;
		X_Re[904] = 15'd35868;
		X_Re[905] = -15'd93185;
		X_Re[906] = -15'd14034;
		X_Re[907] = 15'd24008;
		X_Re[908] = 15'd7848;
		X_Re[909] = 15'd3472;
		X_Re[910] = 15'd8206;
		X_Re[911] = 15'd4331;
		X_Re[912] = -15'd4449;
		X_Re[913] = 15'd7264;
		X_Re[914] = -15'd870;
		X_Re[915] = 15'd13462;
		X_Re[916] = 15'd2968;
		X_Re[917] = 15'd20766;
		X_Re[918] = 15'd36890;
		X_Re[919] = -15'd33732;
		X_Re[920] = -15'd8783;
		X_Re[921] = -15'd6999;
		X_Re[922] = -15'd429;
		X_Re[923] = 15'd2850;
		X_Re[924] = 15'd2743;
		X_Re[925] = 15'd3784;
		X_Re[926] = -15'd6194;
		X_Re[927] = -15'd15483;
		X_Re[928] = -15'd1423;
		X_Re[929] = -15'd32083;
		X_Re[930] = 15'd53368;
		X_Re[931] = 15'd11635;
		X_Re[932] = 15'd10361;
		X_Re[933] = 15'd19519;
		X_Re[934] = 15'd13322;
		X_Re[935] = 15'd328;
		X_Re[936] = 15'd12647;
		X_Re[937] = 15'd6553;
		X_Re[938] = 15'd508;
		X_Re[939] = 15'd1599;
		X_Re[940] = 15'd7487;
		X_Re[941] = 15'd10478;
		X_Re[942] = 15'd5014;
		X_Re[943] = 15'd21865;
		X_Re[944] = -15'd103143;
		X_Re[945] = -15'd322659;
		X_Re[946] = -15'd2159;
		X_Re[947] = 15'd18835;
		X_Re[948] = 15'd15514;
		X_Re[949] = 15'd20953;
		X_Re[950] = 15'd24094;
		X_Re[951] = 15'd27560;
		X_Re[952] = 15'd20529;
		X_Re[953] = 15'd86424;
		X_Re[954] = 15'd24689;
		X_Re[955] = 15'd98286;
		X_Re[956] = 15'd25897;
		X_Re[957] = -15'd220475;
		X_Re[958] = -15'd350559;
		X_Re[959] = -15'd84078;
		X_Re[960] = -15'd89550;
		X_Re[961] = -15'd73725;
		X_Re[962] = -15'd68355;
		X_Re[963] = -15'd76563;
		X_Re[964] = -15'd374488;
		X_Re[965] = 15'd172680;
		X_Re[966] = 15'd99801;
		X_Re[967] = 15'd16164;
		X_Re[968] = 15'd19028;
		X_Re[969] = -15'd2465;
		X_Re[970] = -15'd32042;
		X_Re[971] = 15'd200812;
		X_Re[972] = 15'd3041;
		X_Re[973] = 15'd44296;
		X_Re[974] = 15'd18707;
		X_Re[975] = 15'd19509;
		X_Re[976] = 15'd37484;
		X_Re[977] = 15'd35091;
		X_Re[978] = 15'd7926;
		X_Re[979] = 15'd32371;
		X_Re[980] = 15'd71278;
		X_Re[981] = 15'd19080;
		X_Re[982] = 15'd48085;
		X_Re[983] = 15'd77266;
		X_Re[984] = 15'd422815;
		X_Re[985] = -15'd219111;
		X_Re[986] = -15'd92155;
		X_Re[987] = -15'd33674;
		X_Re[988] = -15'd57943;
		X_Re[989] = 15'd31774;
		X_Re[990] = -15'd22086;
		X_Re[991] = -15'd10798;
		X_Re[992] = -15'd20014;
		X_Re[993] = -15'd23713;
		X_Re[994] = -15'd38433;
		X_Re[995] = -15'd23890;
		X_Re[996] = -15'd34797;
		X_Re[997] = -15'd73347;
		X_Re[998] = 15'd41646;
		X_Re[999] = 15'd2592;
		X_Re[1000] = -15'd5577;
		X_Re[1001] = 15'd13800;
		X_Re[1002] = -15'd4748;
		X_Re[1003] = -15'd19342;
		X_Re[1004] = 15'd1037;
		X_Re[1005] = -15'd54871;
		X_Re[1006] = -15'd32079;
		X_Re[1007] = 15'd41019;
		X_Re[1008] = -15'd12426;
		X_Re[1009] = 15'd16013;
		X_Re[1010] = 15'd2080;
		X_Re[1011] = -15'd40016;
		X_Re[1012] = -15'd7187;
		X_Re[1013] = 15'd71943;
		X_Re[1014] = -15'd45666;
		X_Re[1015] = -15'd166613;
		X_Re[1016] = -15'd5662;
		X_Re[1017] = -15'd45742;
		X_Re[1018] = -15'd13493;
		X_Re[1019] = -15'd8097;
		X_Re[1020] = -15'd3178;
		X_Re[1021] = -15'd3237;
		X_Re[1022] = 15'd8055;
		X_Re[1023] = 15'd3344;	
		#10
		Start = 1;
		//$display("Results 1:");
		//$display("Y[0] expected %d+i%d got %d+i%d", -482739591, 0, Y_Re[0], Y_Im[0]);
		//$display("Y[1] expected %d+i%d got %d+i%d", 322112716, 107370905, Y_Re[1], Y_Im[1]);
		//$display("Y[2] expected %d+i%d got %d+i%d", -161485842, 0, Y_Re[2], Y_Im[2]);
		//$display("Y[3] expected %d+i%d got %d+i%d", 322112716, -107370905, Y_Re[3], Y_Im[3]);
		//#100
		//X_Re[0] = 16'd406;
		//X_Re[1] = 16'd2496;
		//X_Re[2] = 16'd1238;
		//X_Re[3] = -16'd1638;	  
		//#50
		//$display("Results 2:");
		//$display("Y[0] expected %d+i%d got %d+i%d", 164062743, 0, Y_Re[0], Y_Im[0]);
		//$display("Y[1] expected %d+i%d got %d+i%d", -054544420, 271004165, Y_Re[1], Y_Im[1]);
		//$display("Y[2] expected %d+i%d got %d+i%d", 051538034, 0, Y_Re[2], Y_Im[2]);
		//$display("Y[3] expected %d+i%d got %d+i%d", -054544420, -271004165, Y_Re[3], Y_Im[3]);
	end

endmodule